** sch_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/comp_tb-tran.sch
**.subckt comp_tb-tran
VIN in GND PULSE(0V 1.8V 0.5ns 0.1ns 0.1ns 50ns 100ns)
VDD vd GND 1.8
X1 vd out in GND comp
**** begin user architecture code

*cmd step stop
.tran 0.005n 100n
.control
set color0=white
set color1=black
destroy all
run
plot out in 0.9 xlimit 50.45n 50.90n
plot out in

.endc

 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/comp.sym # of pins=4
** sym_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/comp.sym
** sch_path: /home/hugodg/projects-sky130/temp-sensor/sigma-delta_modulator/xschem/comp.sch
.subckt comp  vd out in gnd
*.ipin in
*.iopin gnd
*.opin out
*.iopin vd
**** begin user architecture code




**** end user architecture code
XN1 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XP1 out in vd vd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
