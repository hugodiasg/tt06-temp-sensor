** sch_path: /home/hugodg/projects-sky130/temp-sensor/sensor/xschem/gm-id_1v8.sch
**.subckt gm-id_1v8
VDD vd GND 1.8
Vin vi GND 1.8
XM1 vd vi GND GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.dc vdd 0.1 1.8 0.001
.control
run
set color0=white
set color1=black

let idd=-i(vdd)
let gm_id=1/(abs(vi-vd))

plot idd vs gm_id
.endc



.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
