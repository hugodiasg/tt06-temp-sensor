* NGSPICE file created from sigma-delta_flat.ext - technology: sky130A

.subckt sigma-delta_flat gnd clk out_sigma vts ib out_buff vd out vpwr
X0 gnd.t86 a_15881_829# a_15815_855# gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 vpwr.t3 a_15706_855# a_15881_829# vpwr.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 gnd.t33 gnd.t30 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=1
X3 a_15815_855# a_14625_855# a_15706_855# gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4 a_15046_855# sigma-delta_0.x1.D vpwr.t25 vpwr.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_16688_5320# a_16854_3988# gnd.t120 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X6 buffer_0.a.t15 buffer_0.a.t13 buffer_0.a.t14 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0 ps=0 w=1.5 l=0.15
X7 sensor_0.a.t11 sensor_0.b.t20 gnd.t105 gnd.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X8 sensor_0.b.t15 sensor_0.b.t14 gnd.t106 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X9 a_15430_3152# a_15596_2320# gnd.t91 sky130_fd_pr__res_xhigh_po_0p35 l=2
X10 vd.t15 buffer_0.b.t16 out_buff.t1 vd.t14 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X11 a_14791_855# a_14625_855# gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_15546_5320# sigma-delta_0.in_int gnd.t119 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X13 vd.t43 buffer_0.a.t7 buffer_0.a.t8 vd.t42 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 a_15046_855# sigma-delta_0.x1.D gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X15 gnd.t108 sensor_0.b.t21 vtd.t23 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X16 sensor_0.c sensor_0.c sensor_0.c vd.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=1
X17 buffer_0.d.t4 buffer_0.d.t2 buffer_0.d.t3 vd.t52 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0 w=15 l=1
X18 a_15403_855# a_15359_1097# a_15237_855# gnd.t36 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X19 sigma-delta_0.in_int a_14600_2320# gnd.t75 sky130_fd_pr__res_xhigh_po_0p35 l=2
X20 gnd.t111 ib.t0 ib.t1 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 gnd.t29 gnd.t27 gnd.t28 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X22 a_14550_5320# a_14716_3988# gnd.t132 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X23 ib.t4 ib.t2 ib.t3 gnd.t109 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X24 vpwr.t1 a_15359_1097# a_15249_1221# vpwr.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X25 vts.t16 vtd.t0 vtd.t1 vts.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 gnd.t47 sensor_0.b.t12 sensor_0.b.t13 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X27 a_16356_5320# a_16522_3988# gnd.t44 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X28 gnd.t123 clk.t0 a_14625_855# gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 vtd.t9 vtd.t8 vts.t14 vts.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 gnd.t26 gnd.t24 gnd.t25 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X31 a_15098_3152# a_15264_2320# gnd.t90 sky130_fd_pr__res_xhigh_po_0p35 l=2
X32 vpwr.t5 clk.t1 a_14625_855# vpwr.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X33 gnd.t131 sensor_0.b.t22 sensor_0.a.t10 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X34 gnd.t23 gnd.t21 gnd.t22 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X35 vtd.t22 sensor_0.b.t23 gnd.t133 gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X36 vts.t12 vtd.t14 vtd.t15 vts.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 buffer_0.b.t12 buffer_0.b.t11 vd.t13 vd.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X38 gnd.t74 sigma-delta_0.in_comp sigma-delta_0.x1.D gnd.t73 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X39 vtd.t21 sensor_0.b.t24 gnd.t134 gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X40 a_17020_5320# sigma-delta_0.x1.Q gnd.t35 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X41 vtd.t11 vtd.t10 vts.t10 vts.t9 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X42 vd.t11 buffer_0.b.t5 buffer_0.b.t6 vd.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X43 sigma-delta_0.x1.Q a_15881_829# vpwr.t23 vpwr.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.213 ps=1.67 w=1 l=0.15
X44 a_15359_1097# a_15141_855# gnd.t113 gnd.t112 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X45 vd.t53 a_6126_29386# gnd.t118 sky130_fd_pr__res_xhigh_po_0p35 l=5
X46 sensor_0.b.t17 vtd.t24 sensor_0.c vd.t47 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X47 sigma-delta_0.in_comp gnd.t72 sky130_fd_pr__cap_mim_m3_2 l=27.2 w=27.2
X48 a_16060_855# vpwr.t30 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X49 vts.t8 vtd.t2 vtd.t3 vts.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X50 vd.t9 buffer_0.b.t9 buffer_0.b.t10 vd.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X51 gnd.t107 sensor_0.b.t10 sensor_0.b.t11 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X52 buffer_0.a.t12 buffer_0.a.t11 buffer_0.a.t12 vd.t41 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X53 vd.t26 sensor_0.a.t0 sensor_0.a.t1 vd.t25 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X54 buffer_0.a.t4 buffer_0.a.t3 vd.t40 vd.t39 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X55 buffer_0.b.t15 vts.t25 buffer_0.c gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X56 sensor_0.b.t9 sensor_0.b.t8 gnd.t66 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X57 a_14882_5320# a_15048_3988# gnd.t137 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X58 gnd.t101 sensor_0.b.t25 sensor_0.a.t9 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X59 vpwr.t21 a_15881_829# a_15868_1221# vpwr.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X60 a_15881_829# a_15706_855# a_16060_855# gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X61 vts.t24 vts.t21 vts.t23 vts.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X62 buffer_0.d.t11 buffer_0.a.t16 vd.t38 vd.t37 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X63 out_buff.t10 buffer_0.d.t9 sky130_fd_pr__cap_mim_m3_2 l=15 w=30
X64 gnd.t129 sensor_0.b.t26 vtd.t20 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X65 vd.t51 vtd.t25 vts.t6 vd.t50 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
X66 a_15214_5320# a_15380_3988# gnd.t136 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X67 vd.t72 vd.t69 vd.t71 vd.t70 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X68 gnd.t20 gnd.t18 gnd.t19 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X69 sensor_0.c vtd.t26 sensor_0.b.t16 vd.t46 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X70 out_buff.t9 out_buff.t7 out_buff.t8 vd.t28 sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=0 ps=0 w=15 l=1
X71 sigma-delta_0.in_comp a_15596_2320# gnd.t127 sky130_fd_pr__res_xhigh_po_0p35 l=2
X72 vd.t68 vd.t65 vd.t67 vd.t66 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X73 sensor_0.a.t8 sensor_0.b.t27 gnd.t128 gnd.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X74 sensor_0.a.t7 sensor_0.b.t28 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X75 sensor_0.a.t3 sensor_0.a.t2 vd.t24 vd.t23 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X76 gnd.t68 buffer_0.d.t12 out_buff.t3 gnd.t67 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X77 vd.t73 out.t3 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X78 a_14766_3152# a_14600_2320# gnd.t98 sky130_fd_pr__res_xhigh_po_0p35 l=2
X79 buffer_0.c out_buff.t11 buffer_0.a.t0 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X80 out_buff.t2 buffer_0.d.t13 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_16024_5320# a_16190_3988# gnd.t126 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X82 sensor_0.b.t7 sensor_0.b.t6 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X83 vd.t64 vd.t62 vd.t64 vd.t63 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=1
X84 gnd.t125 buffer_0.d.t7 buffer_0.d.t8 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 gnd.t43 sensor_0.b.t29 vtd.t19 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X86 a_15249_1221# a_14625_855# a_15141_855# vpwr.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X87 a_16688_5320# a_16522_3988# gnd.t103 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X88 vd.t61 vd.t58 vd.t60 vd.t59 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X89 vd.t7 buffer_0.b.t7 buffer_0.b.t8 vd.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X90 buffer_0.d.t6 buffer_0.d.t5 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 sensor_0.c sensor_0.a.t12 sensor_0.d vd.t22 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X92 a_15430_3152# a_15264_2320# gnd.t89 sky130_fd_pr__res_xhigh_po_0p35 l=2
X93 sensor_0.d sensor_0.a.t13 sensor_0.c vd.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X94 a_15546_5320# a_15380_3988# gnd.t60 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X95 buffer_0.d.t1 buffer_0.d.t0 buffer_0.d.t1 vd.t0 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0 w=15 l=1
X96 gnd.t17 gnd.t15 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=1
X97 gnd.t14 gnd.t12 gnd.t13 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X98 gnd.t11 gnd.t9 gnd.t10 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X99 a_15249_1221# vpwr.t11 vpwr.t13 vpwr.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X100 gnd.t8 gnd.t5 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X101 buffer_0.c buffer_0.c buffer_0.c gnd.t63 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=1.08 ps=8.82 w=1 l=1
X102 vd.t57 vd.t54 vd.t56 vd.t55 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X103 a_15881_829# vpwr.t8 vpwr.t10 vpwr.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X104 vtd.t5 vtd.t4 vts.t5 vts.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X105 vd.t36 buffer_0.a.t17 buffer_0.d.t10 vd.t35 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X106 sigma-delta_0.in_int gnd.t76 sky130_fd_pr__cap_mim_m3_2 l=27.2 w=27.2
X107 gnd.t41 sensor_0.b.t4 sensor_0.b.t5 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X108 buffer_0.c ib.t5 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X109 vts.t3 vtd.t12 vtd.t13 vts.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X110 buffer_0.b.t4 buffer_0.b.t2 buffer_0.b.t3 vd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X111 vd.t17 sigma-delta_0.in_comp sigma-delta_0.x1.D vd.t16 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X112 gnd.t102 sensor_0.b.t30 sensor_0.a.t6 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X113 vtd.t18 sensor_0.b.t31 gnd.t71 gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X114 a_16356_5320# a_16190_3988# gnd.t0 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X115 vtd.t7 vtd.t6 vts.t1 vts.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X116 sigma-delta_0.x1.Q a_15881_829# gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X117 vtd.t17 sensor_0.b.t32 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X118 a_15098_3152# a_14932_2320# gnd.t95 sky130_fd_pr__res_xhigh_po_0p35 l=2
X119 a_15706_855# a_14791_855# a_15359_1097# gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X120 sensor_0.c vtd.t27 sensor_0.b.t19 vd.t49 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X121 out_buff.t0 buffer_0.b.t17 vd.t4 vd.t3 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X122 a_15214_5320# a_15048_3988# gnd.t53 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X123 buffer_0.a.t10 buffer_0.a.t9 vd.t34 vd.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X124 vd.t74 out.t2 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X125 gnd.t82 a_15881_829# a_16445_855# gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X126 a_15868_1221# a_14791_855# a_15706_855# vpwr.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X127 a_14791_855# a_14625_855# vpwr.t16 vpwr.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X128 vd.t32 buffer_0.a.t1 buffer_0.a.t2 vd.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X129 sensor_0.b.t18 vtd.t28 sensor_0.c vd.t48 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X130 a_17020_5320# a_16854_3988# gnd.t34 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X131 gnd.t69 sensor_0.b.t2 sensor_0.b.t3 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X132 sensor_0.d vtd.t29 vd.t45 vd.t44 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X133 buffer_0.a.t6 buffer_0.a.t5 vd.t30 vd.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X134 a_14882_5320# a_14716_3988# gnd.t115 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X135 a_15141_855# a_14791_855# a_15046_855# vpwr.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X136 sensor_0.d sensor_0.a.t14 sensor_0.c vd.t20 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X137 vts.t20 vts.t17 vts.t19 vts.t18 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X138 buffer_0.b.t1 buffer_0.b.t0 buffer_0.b.t1 gnd.t114 sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0 ps=0 w=1.5 l=0.15
X139 sensor_0.b.t1 sensor_0.b.t0 gnd.t135 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X140 gnd.t100 sensor_0.b.t33 sensor_0.a.t5 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X141 a_16024_5320# sigma-delta_0.in_int gnd.t121 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X142 vd.t75 out.t1 sky130_fd_pr__cap_mim_m3_2 l=24.4 w=24.4
X143 a_15141_855# a_14625_855# a_15046_855# gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X144 gnd.t52 out_sigma.t2 out.t0 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X145 sensor_0.c sensor_0.a.t15 sensor_0.d vd.t19 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X146 gnd.t104 sensor_0.b.t34 vtd.t16 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X147 a_15237_855# a_14791_855# a_15141_855# gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X148 out_sigma.t1 a_16445_855# vpwr.t29 vpwr.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X149 vpwr.t19 a_15881_829# a_16445_855# vpwr.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X150 gnd.t58 vpwr.t31 a_15403_855# gnd.t57 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X151 out_sigma.t0 a_16445_855# gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X152 a_15706_855# a_14625_855# a_15359_1097# vpwr.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X153 a_14550_5320# out_buff.t4 gnd.t70 sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X154 sensor_0.a.t4 sensor_0.b.t35 gnd.t54 gnd.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X155 a_14766_3152# a_14932_2320# gnd.t59 sky130_fd_pr__res_xhigh_po_0p35 l=2
X156 a_15359_1097# a_15141_855# vpwr.t27 vpwr.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X157 gnd.t4 gnd.t1 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X158 buffer_0.b.t14 buffer_0.b.t13 vd.t2 vd.t1 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X159 out_buff.t6 out_buff.t5 out_buff.t6 vd.t27 sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=0 ps=0 w=15 l=1
R0 gnd.n164 gnd.n3 16393.5
R1 gnd.n149 gnd.n143 9351.88
R2 gnd.n162 gnd.n11 7246.65
R3 gnd.n164 gnd.n163 4031.02
R4 gnd.n163 gnd.n162 2559.7
R5 gnd.n161 gnd 1652.19
R6 gnd.n142 gnd.n136 1498.93
R7 gnd.n140 gnd.n139 1273.6
R8 gnd.n9 gnd.n8 1273.6
R9 gnd.n162 gnd.n161 1184.7
R10 gnd.n167 gnd.n164 1057.91
R11 gnd.n143 gnd.n142 759.644
R12 gnd.n205 gnd.n204 585
R13 gnd.n259 gnd.n258 585
R14 gnd.n261 gnd.n260 585
R15 gnd.n2 gnd.n1 585
R16 gnd.n30 gnd.n27 560.566
R17 gnd.n38 gnd.n35 547.013
R18 gnd.n131 gnd.n130 523.47
R19 gnd.n28 gnd.t16 348.421
R20 gnd.n137 gnd.t35 342.634
R21 gnd.n169 gnd.t55 334.93
R22 gnd.n267 gnd.t99 331.329
R23 gnd.t116 gnd.n160 330.392
R24 gnd.t78 gnd.t92 307.483
R25 gnd.t114 gnd.t96 305.267
R26 gnd.t40 gnd.n206 298.916
R27 gnd.t130 gnd.t63 263.712
R28 gnd.n207 gnd.t64 262.902
R29 gnd.n43 gnd.n41 256.471
R30 gnd.n130 gnd.n129 247.828
R31 gnd.n51 gnd.n48 242.918
R32 gnd.t83 gnd.t81 226.692
R33 gnd.t37 gnd.t83 226.692
R34 gnd.n160 gnd.n159 224.325
R35 gnd.n235 gnd.t42 223.286
R36 gnd.n49 gnd.t124 217.363
R37 gnd.n59 gnd.t93 215.036
R38 gnd.n39 gnd.t110 214.167
R39 gnd.t35 gnd.t34 204.595
R40 gnd.t103 gnd.t120 204.595
R41 gnd.t44 gnd.t103 204.595
R42 gnd.t0 gnd.t44 204.595
R43 gnd.t126 gnd.t0 204.595
R44 gnd.t121 gnd.t126 204.595
R45 gnd.t49 gnd.t36 200.165
R46 gnd.n39 gnd.t87 198.185
R47 gnd.n6 gnd.t127 195.966
R48 gnd.n49 gnd.t61 194.988
R49 gnd.t85 gnd.t45 179.667
R50 gnd.t6 gnd.n168 172.868
R51 gnd.n237 gnd.n234 163.766
R52 gnd.t57 gnd.t112 159.167
R53 gnd.n269 gnd.n259 156.236
R54 gnd.n69 gnd.t84 154.317
R55 gnd.n216 gnd.n215 153.976
R56 gnd.t48 gnd.t130 153.434
R57 gnd.n168 gnd.n167 152.16
R58 gnd.n214 gnd.n209 150.648
R59 gnd.n157 gnd.n156 149.835
R60 gnd.n216 gnd.n205 148.707
R61 gnd.n51 gnd.n30 147.294
R62 gnd.t89 gnd.t60 142.97
R63 gnd.t90 gnd.t136 142.97
R64 gnd.t95 gnd.t53 142.97
R65 gnd.t59 gnd.t137 142.97
R66 gnd.t98 gnd.t115 142.97
R67 gnd.t75 gnd.t132 142.97
R68 gnd.n41 gnd.n38 133.742
R69 gnd.t50 gnd.t80 131.434
R70 gnd.n71 gnd.n70 128.757
R71 gnd.t2 gnd.n266 127.85
R72 gnd.n6 gnd.t121 126.948
R73 gnd.t112 gnd.t50 119.376
R74 gnd.n235 gnd.t38 118.847
R75 gnd.t81 gnd.t116 116.965
R76 gnd.n67 gnd.n66 116.754
R77 gnd.t80 gnd.t85 115.758
R78 gnd.t77 gnd.t49 115.758
R79 gnd.t92 gnd.t77 114.552
R80 gnd.n266 gnd.n265 110.743
R81 gnd.t45 gnd.t37 109.73
R82 gnd.n11 gnd.n5 108.46
R83 gnd.n98 gnd.n57 107.24
R84 gnd.n85 gnd.n63 107.24
R85 gnd.t31 gnd.t114 107.084
R86 gnd.n5 gnd.t70 103.529
R87 gnd.t122 gnd.t78 101.288
R88 gnd.n66 gnd.t46 100.001
R89 gnd.n156 gnd.n152 98.6358
R90 gnd.t36 gnd.t57 86.8188
R91 gnd.n163 gnd.n4 86.3064
R92 gnd.n207 gnd.t40 79.2311
R93 gnd gnd.t122 78.3781
R94 gnd.n63 gnd.t58 72.8576
R95 gnd.n66 gnd.t86 70.0005
R96 gnd.n171 gnd.n2 65.8829
R97 gnd.n21 gnd.t30 65.675
R98 gnd.n15 gnd.t15 65.5414
R99 gnd.t99 gnd.n262 64.8256
R100 gnd.n28 gnd.t67 63.9308
R101 gnd.t127 gnd.t119 61.6251
R102 gnd.t60 gnd.t91 61.6251
R103 gnd.t136 gnd.t89 61.6251
R104 gnd.t53 gnd.t90 61.6251
R105 gnd.t137 gnd.t95 61.6251
R106 gnd.t115 gnd.t59 61.6251
R107 gnd.t132 gnd.t98 61.6251
R108 gnd.t70 gnd.t75 61.6251
R109 gnd.n63 gnd.t113 60.5809
R110 gnd.n70 gnd.t82 57.1434
R111 gnd.n269 gnd.n261 48.5652
R112 gnd.n57 gnd.t79 38.5719
R113 gnd.n57 gnd.t123 38.5719
R114 gnd.n251 gnd.t1 37.3602
R115 gnd.n254 gnd.t27 37.3602
R116 gnd.n257 gnd.t9 37.3602
R117 gnd.n176 gnd.t21 37.3602
R118 gnd.n179 gnd.t12 37.3602
R119 gnd.n182 gnd.t24 37.3602
R120 gnd.n46 gnd.t31 35.1621
R121 gnd.n87 gnd.n86 34.6358
R122 gnd.n87 gnd.n61 34.6358
R123 gnd.n91 gnd.n61 34.6358
R124 gnd.n92 gnd.n91 34.6358
R125 gnd.n93 gnd.n92 34.6358
R126 gnd.n79 gnd.n78 34.6358
R127 gnd.n80 gnd.n79 34.6358
R128 gnd.n80 gnd.n64 34.6358
R129 gnd.n84 gnd.n64 34.6358
R130 gnd.n74 gnd.n73 34.6358
R131 gnd.n75 gnd.n74 34.6358
R132 gnd.n97 gnd.n59 29.7417
R133 gnd.n73 gnd.n69 27.8593
R134 gnd.n70 gnd.t117 25.4291
R135 gnd.n129 gnd.t51 24.5503
R136 gnd.n99 gnd.n98 24.4919
R137 gnd.n120 gnd.n117 24.3682
R138 gnd.n213 gnd.n210 23.4095
R139 gnd.n136 gnd.t118 22.9965
R140 gnd.t118 gnd.n131 22.9965
R141 gnd.n98 gnd.n97 22.9652
R142 gnd.n163 gnd.t48 20.7778
R143 gnd.n173 gnd.t5 18.6812
R144 gnd.n248 gnd.t18 18.6809
R145 gnd.n75 gnd.n67 17.6946
R146 gnd.n231 gnd.t129 17.4089
R147 gnd.n201 gnd.t69 17.4089
R148 gnd.n242 gnd.t131 17.4084
R149 gnd.n240 gnd.t100 17.4084
R150 gnd.n239 gnd.t101 17.4084
R151 gnd.n242 gnd.t128 17.4084
R152 gnd.n240 gnd.t39 17.4084
R153 gnd.n239 gnd.t54 17.4084
R154 gnd.n231 gnd.t65 17.4079
R155 gnd.n201 gnd.t135 17.4079
R156 gnd.n244 gnd.t105 17.4074
R157 gnd.n244 gnd.t102 17.4074
R158 gnd.n218 gnd.t43 17.4069
R159 gnd.n218 gnd.t133 17.4055
R160 gnd.n247 gnd.t20 17.405
R161 gnd.n247 gnd.t19 17.405
R162 gnd.n250 gnd.t4 17.405
R163 gnd.n250 gnd.t3 17.405
R164 gnd.n253 gnd.t29 17.405
R165 gnd.n253 gnd.t28 17.405
R166 gnd.n256 gnd.t11 17.405
R167 gnd.n256 gnd.t10 17.405
R168 gnd.n172 gnd.t8 17.405
R169 gnd.n172 gnd.t7 17.405
R170 gnd.n175 gnd.t23 17.405
R171 gnd.n175 gnd.t22 17.405
R172 gnd.n178 gnd.t14 17.405
R173 gnd.n178 gnd.t13 17.405
R174 gnd.n181 gnd.t26 17.405
R175 gnd.n181 gnd.t25 17.405
R176 gnd.n13 gnd.t74 17.405
R177 gnd.n220 gnd.t71 17.4034
R178 gnd.n219 gnd.t108 17.4034
R179 gnd.n226 gnd.t134 17.4034
R180 gnd.n225 gnd.t104 17.4034
R181 gnd.n196 gnd.t66 17.4034
R182 gnd.n195 gnd.t107 17.4034
R183 gnd.n190 gnd.t56 17.4034
R184 gnd.n189 gnd.t41 17.4034
R185 gnd.n185 gnd.t106 17.4034
R186 gnd.n184 gnd.t47 17.4034
R187 gnd.n31 gnd.t88 17.4005
R188 gnd.n31 gnd.t111 17.4005
R189 gnd.n93 gnd.n59 14.6829
R190 gnd.n48 gnd.n43 13.5534
R191 gnd.n36 gnd.t109 12.7866
R192 gnd.n46 gnd.t94 11.1883
R193 gnd.n71 gnd.n69 10.9075
R194 gnd.n267 gnd.t2 10.8047
R195 gnd.n13 gnd.n12 9.33321
R196 gnd.n171 gnd.n170 9.3005
R197 gnd.n170 gnd.n169 9.3005
R198 gnd.n216 gnd.n208 9.3005
R199 gnd.n208 gnd.n207 9.3005
R200 gnd.n237 gnd.n236 9.3005
R201 gnd.n236 gnd.n235 9.3005
R202 gnd.n269 gnd.n268 9.3005
R203 gnd.n268 gnd.n267 9.3005
R204 gnd.n125 gnd.t52 8.70236
R205 gnd.n86 gnd.n85 7.90638
R206 gnd.n169 gnd.t6 7.20328
R207 gnd.n21 gnd.t33 6.44128
R208 gnd.n53 gnd.n52 5.41306
R209 gnd.n33 gnd.n32 5.41306
R210 gnd.n95 gnd.n59 4.6505
R211 gnd.n73 gnd.n72 4.6505
R212 gnd.n74 gnd.n68 4.6505
R213 gnd.n76 gnd.n75 4.6505
R214 gnd.n78 gnd.n77 4.6505
R215 gnd.n79 gnd.n65 4.6505
R216 gnd.n81 gnd.n80 4.6505
R217 gnd.n82 gnd.n64 4.6505
R218 gnd.n84 gnd.n83 4.6505
R219 gnd.n86 gnd.n62 4.6505
R220 gnd.n88 gnd.n87 4.6505
R221 gnd.n89 gnd.n61 4.6505
R222 gnd.n91 gnd.n90 4.6505
R223 gnd.n92 gnd.n60 4.6505
R224 gnd.n94 gnd.n93 4.6505
R225 gnd.n97 gnd.n96 4.6505
R226 gnd.n98 gnd.n58 4.6505
R227 gnd.n55 gnd.n54 4.5005
R228 gnd.n56 gnd.n54 4.5005
R229 gnd.n18 gnd.t62 3.4805
R230 gnd.n18 gnd.t125 3.4805
R231 gnd.n16 gnd.t17 3.4805
R232 gnd.n16 gnd.t68 3.4805
R233 gnd.n22 gnd.t97 3.4805
R234 gnd.n22 gnd.t32 3.4805
R235 gnd.n17 gnd.n15 3.21916
R236 gnd.n23 gnd.n21 2.95318
R237 gnd.n78 gnd.n67 2.63579
R238 gnd.n125 gnd 2.5773
R239 gnd.n103 gnd.n53 2.43634
R240 gnd.n100 gnd.n54 2.25328
R241 gnd gnd.n0 2.00418
R242 gnd.n104 gnd.n14 1.93469
R243 gnd.n85 gnd.n84 1.88285
R244 gnd gnd.n102 1.72422
R245 gnd.n33 gnd.n31 1.41862
R246 gnd.n104 gnd.n103 1.22706
R247 gnd gnd.n0 1.2022
R248 gnd.n32 gnd 0.793114
R249 gnd.n273 gnd.n272 0.685777
R250 gnd.n20 gnd.n17 0.6455
R251 gnd.n24 gnd.n23 0.62925
R252 gnd.n106 gnd.n104 0.575502
R253 gnd.n151 gnd.n150 0.54125
R254 gnd.n152 gnd.n151 0.541165
R255 gnd.n224 gnd.n218 0.447415
R256 gnd.n230 gnd.n224 0.438
R257 gnd.n232 gnd.n230 0.438
R258 gnd.n52 gnd.n25 0.425505
R259 gnd.n194 gnd.n188 0.375501
R260 gnd.n233 gnd.n232 0.375501
R261 gnd.n200 gnd.n194 0.3755
R262 gnd.n202 gnd.n200 0.3755
R263 gnd.n241 gnd.n239 0.373217
R264 gnd.n243 gnd.n241 0.371401
R265 gnd.n245 gnd.n243 0.369555
R266 gnd.n128 gnd.n124 0.366293
R267 gnd.n115 gnd.n114 0.365897
R268 gnd.n129 gnd.n115 0.365897
R269 gnd.n124 gnd.n123 0.365897
R270 gnd.n148 gnd.n147 0.347558
R271 gnd.n147 gnd.n146 0.347269
R272 gnd.n246 gnd.n245 0.338503
R273 gnd.n203 gnd.n202 0.330858
R274 gnd.n203 gnd.n183 0.290469
R275 gnd.n233 gnd.n217 0.281539
R276 gnd.n14 gnd.t72 0.266467
R277 gnd.n238 gnd.n233 0.245825
R278 gnd.n271 gnd.n246 0.244548
R279 gnd.n273 gnd.n0 0.230614
R280 gnd.n246 gnd.n238 0.180349
R281 gnd.n217 gnd.n203 0.156539
R282 gnd.n72 gnd.n71 0.144332
R283 gnd.n111 gnd.n110 0.1305
R284 gnd.t118 gnd.n111 0.1305
R285 gnd.n133 gnd.n132 0.1305
R286 gnd.t118 gnd.n133 0.1305
R287 gnd.n72 gnd.n68 0.120292
R288 gnd.n76 gnd.n68 0.120292
R289 gnd.n77 gnd.n76 0.120292
R290 gnd.n77 gnd.n65 0.120292
R291 gnd.n81 gnd.n65 0.120292
R292 gnd.n82 gnd.n81 0.120292
R293 gnd.n83 gnd.n82 0.120292
R294 gnd.n83 gnd.n62 0.120292
R295 gnd.n88 gnd.n62 0.120292
R296 gnd.n89 gnd.n88 0.120292
R297 gnd.n90 gnd.n89 0.120292
R298 gnd.n90 gnd.n60 0.120292
R299 gnd.n94 gnd.n60 0.120292
R300 gnd.n95 gnd.n94 0.120292
R301 gnd.n96 gnd.n95 0.120292
R302 gnd.n96 gnd.n58 0.120292
R303 gnd.n154 gnd.n153 0.10956
R304 gnd.t73 gnd.n154 0.10956
R305 gnd.n155 gnd.t73 0.10956
R306 gnd.n156 gnd.n155 0.10956
R307 gnd.n119 gnd.n118 0.10956
R308 gnd.n122 gnd.n121 0.10956
R309 gnd.t51 gnd.n122 0.10956
R310 gnd.n120 gnd.n119 0.109135
R311 gnd.n148 gnd.n145 0.0849523
R312 gnd.n145 gnd.n144 0.0845034
R313 gnd.n274 gnd.n273 0.0772045
R314 gnd.n274 gnd 0.0755
R315 gnd.n58 gnd.n55 0.0734167
R316 gnd.n249 gnd.n248 0.073412
R317 gnd.n174 gnd.n173 0.0734113
R318 gnd.n25 gnd.n24 0.063
R319 gnd.n175 gnd.n174 0.0610469
R320 gnd.n176 gnd.n175 0.0610469
R321 gnd.n178 gnd.n177 0.0610469
R322 gnd.n179 gnd.n178 0.0610469
R323 gnd.n181 gnd.n180 0.0610469
R324 gnd.n182 gnd.n181 0.0610469
R325 gnd.n250 gnd.n249 0.0610469
R326 gnd.n251 gnd.n250 0.0610469
R327 gnd.n253 gnd.n252 0.0610469
R328 gnd.n254 gnd.n253 0.0610469
R329 gnd.n256 gnd.n255 0.0610469
R330 gnd.n257 gnd.n256 0.0610469
R331 gnd.n270 gnd.n257 0.0573558
R332 gnd.n183 gnd.n182 0.0573547
R333 gnd.n271 gnd.n270 0.0464211
R334 gnd.n38 gnd.n37 0.0431634
R335 gnd.n37 gnd.n36 0.0431634
R336 gnd.n177 gnd.n176 0.0426875
R337 gnd.n180 gnd.n179 0.0426875
R338 gnd.n252 gnd.n251 0.0426875
R339 gnd.n255 gnd.n254 0.0426875
R340 gnd.n158 gnd.n157 0.0425017
R341 gnd.n159 gnd.n158 0.0425017
R342 gnd.n272 gnd 0.0395625
R343 gnd.n30 gnd.n29 0.0388129
R344 gnd.n29 gnd.n28 0.0388129
R345 gnd gnd.n274 0.0345909
R346 gnd.n56 gnd 0.0330521
R347 gnd.n103 gnd 0.03175
R348 gnd.n173 gnd.n172 0.031274
R349 gnd.n248 gnd.n247 0.0312734
R350 gnd.n101 gnd.n55 0.0265417
R351 gnd.n117 gnd.n116 0.0264102
R352 gnd.n99 gnd 0.0226354
R353 gnd.n43 gnd.n42 0.0215341
R354 gnd.n42 gnd.n4 0.0215341
R355 gnd.n24 gnd.n20 0.01675
R356 gnd.n232 gnd.n231 0.0153409
R357 gnd.n229 gnd.n227 0.0129048
R358 gnd.n101 gnd.n100 0.0114272
R359 gnd.n223 gnd.n221 0.0114167
R360 gnd.n100 gnd.n99 0.0113582
R361 gnd.n102 gnd.n54 0.0110001
R362 gnd.n48 gnd.n47 0.00984699
R363 gnd.n47 gnd.n46 0.00984699
R364 gnd.n215 gnd.n214 0.0092427
R365 gnd.n214 gnd.n213 0.0092427
R366 gnd.n264 gnd.n263 0.00883856
R367 gnd.n265 gnd.n264 0.00883856
R368 gnd.n166 gnd.n165 0.00883856
R369 gnd.n167 gnd.n166 0.00883856
R370 gnd.n107 gnd.n13 0.00867757
R371 gnd.n202 gnd.n201 0.00792873
R372 gnd.n113 gnd.n112 0.00762598
R373 gnd.n131 gnd.n113 0.00762598
R374 gnd.n135 gnd.n134 0.00762598
R375 gnd.n136 gnd.n135 0.00762598
R376 gnd.n27 gnd.n26 0.007537
R377 gnd.n35 gnd.n34 0.007537
R378 gnd.n41 gnd.n40 0.00701261
R379 gnd.n40 gnd.n39 0.00701261
R380 gnd.n51 gnd.n50 0.00701261
R381 gnd.n50 gnd.n49 0.00701261
R382 gnd.n107 gnd.n106 0.00634112
R383 gnd gnd.n56 0.00570833
R384 gnd.n199 gnd.n197 0.00546432
R385 gnd.n45 gnd.n44 0.00517349
R386 gnd.n46 gnd.n45 0.00517349
R387 gnd.n8 gnd.n7 0.00517349
R388 gnd.n7 gnd.n6 0.00517349
R389 gnd.n141 gnd.n140 0.00517349
R390 gnd.n142 gnd.n141 0.00517349
R391 gnd.n186 gnd.n184 0.00502806
R392 gnd.n191 gnd.n189 0.00502806
R393 gnd.n197 gnd.n195 0.00502805
R394 gnd.n221 gnd.n219 0.00502803
R395 gnd.n227 gnd.n225 0.00502803
R396 gnd.n212 gnd.n211 0.00487141
R397 gnd.n213 gnd.n212 0.00487141
R398 gnd.n150 gnd.n109 0.00441022
R399 gnd.n10 gnd.n9 0.0043402
R400 gnd.n11 gnd.n10 0.0043402
R401 gnd.n139 gnd.n138 0.0043402
R402 gnd.n138 gnd.n137 0.0043402
R403 gnd.n186 gnd.n185 0.00402807
R404 gnd.n191 gnd.n190 0.00402806
R405 gnd.n197 gnd.n196 0.00402806
R406 gnd.n221 gnd.n220 0.00402804
R407 gnd.n227 gnd.n226 0.00402803
R408 gnd.n193 gnd.n191 0.00397623
R409 gnd.n109 gnd.n108 0.00391284
R410 gnd.n108 gnd.n107 0.00391159
R411 gnd.n20 gnd.n19 0.00371923
R412 gnd.n17 gnd.n16 0.00294771
R413 gnd.n23 gnd.n22 0.00294771
R414 gnd.n14 gnd.t76 0.00288363
R415 gnd.n188 gnd.n186 0.00248813
R416 gnd.n272 gnd.n271 0.00245312
R417 gnd.n128 gnd.n127 0.00236777
R418 gnd.n19 gnd.n18 0.00217489
R419 gnd.t51 gnd.n120 0.00192099
R420 gnd.n127 gnd.n126 0.00186816
R421 gnd.n270 gnd.n269 0.00152216
R422 gnd.n183 gnd.n171 0.00152195
R423 gnd.n41 gnd.n33 0.00148887
R424 gnd.n52 gnd.n51 0.00148887
R425 gnd.n229 gnd.n228 0.00138337
R426 gnd.n223 gnd.n222 0.00138109
R427 gnd.n199 gnd.n198 0.00134613
R428 gnd.n193 gnd.n192 0.00134049
R429 gnd.n188 gnd.n187 0.001335
R430 gnd.n126 gnd.n125 0.00124275
R431 gnd.n243 gnd.n242 0.00121065
R432 gnd.n241 gnd.n240 0.001204
R433 gnd.n149 gnd.n148 0.00104118
R434 gnd.n102 gnd.n101 0.00100955
R435 gnd.n150 gnd.n149 0.00100261
R436 gnd.n245 gnd.n244 0.00100079
R437 gnd.n129 gnd.n128 0.00100039
R438 gnd.n217 gnd.n216 0.000522345
R439 gnd.n238 gnd.n237 0.000522345
R440 gnd.n106 gnd.n105 0.00051897
R441 gnd.n230 gnd.n229 0.000501021
R442 gnd.n224 gnd.n223 0.000501021
R443 gnd.n194 gnd.n193 0.000500672
R444 gnd.n200 gnd.n199 0.000500672
R445 vpwr.t15 vpwr.t24 790.188
R446 vpwr.t22 vpwr.t18 648.131
R447 vpwr.t12 vpwr.t26 583.023
R448 vpwr.n77 vpwr 548.548
R449 vpwr.n56 vpwr.t27 514.011
R450 vpwr.t2 vpwr.t22 485.358
R451 vpwr.t17 vpwr.t0 414.33
R452 vpwr.n14 vpwr.t11 413.315
R453 vpwr.n32 vpwr.t25 375.277
R454 vpwr.n7 vpwr.t8 344.005
R455 vpwr.t20 vpwr.t9 319.627
R456 vpwr.n50 vpwr.n39 311.957
R457 vpwr.n72 vpwr.n31 311.894
R458 vpwr.n59 vpwr.n58 309.18
R459 vpwr.t26 vpwr.t14 292.991
R460 vpwr.t6 vpwr.t17 292.991
R461 vpwr.n43 vpwr.n40 292.5
R462 vpwr.n45 vpwr.n44 292.5
R463 vpwr.t18 vpwr.t28 287.072
R464 vpwr.t0 vpwr.t12 287.072
R465 vpwr.t24 vpwr.t6 272.274
R466 vpwr.t14 vpwr.t7 254.518
R467 vpwr.t9 vpwr.t2 248.599
R468 vpwr.t7 vpwr.t20 248.599
R469 vpwr.t4 vpwr.t15 244.306
R470 vpwr.n6 vpwr.t30 187.321
R471 vpwr vpwr.t4 186.556
R472 vpwr.n44 vpwr.n43 182.929
R473 vpwr.n7 vpwr.n5 152
R474 vpwr.n42 vpwr.n41 148.689
R475 vpwr.n14 vpwr.t31 126.127
R476 vpwr.n39 vpwr.t21 119.608
R477 vpwr.n58 vpwr.t1 93.81
R478 vpwr.n6 vpwr.n1 73.2067
R479 vpwr.n43 vpwr.t3 68.0124
R480 vpwr.n58 vpwr.t13 63.3219
R481 vpwr.n39 vpwr.t10 63.3219
R482 vpwr.n41 vpwr.t19 61.9158
R483 vpwr.n31 vpwr.t16 41.5552
R484 vpwr.n31 vpwr.t5 41.5552
R485 vpwr.n71 vpwr.n70 34.6358
R486 vpwr.n64 vpwr.n34 34.6358
R487 vpwr.n65 vpwr.n64 34.6358
R488 vpwr.n66 vpwr.n65 34.6358
R489 vpwr.n60 vpwr.n57 34.6358
R490 vpwr.n51 vpwr.n37 34.6358
R491 vpwr.n55 vpwr.n37 34.6358
R492 vpwr.n66 vpwr.n32 32.377
R493 vpwr.n56 vpwr.n55 32.0005
R494 vpwr.n41 vpwr.t29 30.239
R495 vpwr.n50 vpwr.n49 30.1181
R496 vpwr.n44 vpwr.t23 29.316
R497 vpwr.n72 vpwr.n71 22.9652
R498 vpwr.n51 vpwr.n50 20.3299
R499 vpwr.n70 vpwr.n32 18.0711
R500 vpwr vpwr.n4 14.0185
R501 vpwr.n45 vpwr.n42 13.9946
R502 vpwr.n49 vpwr.n40 12.8758
R503 vpwr.n57 vpwr.n56 9.41227
R504 vpwr.n11 vpwr.n10 9.3005
R505 vpwr.n8 vpwr.n2 9.3005
R506 vpwr.n8 vpwr.n7 9.3005
R507 vpwr.n7 vpwr.n6 9.15991
R508 vpwr.n15 vpwr.n14 7.02651
R509 vpwr.n59 vpwr.n34 6.02403
R510 vpwr.n46 vpwr.n45 5.00414
R511 vpwr.n4 vpwr 4.7293
R512 vpwr.n9 vpwr.n0 4.6505
R513 vpwr.n18 vpwr.n17 4.6505
R514 vpwr.n47 vpwr.n46 4.6505
R515 vpwr.n49 vpwr.n48 4.6505
R516 vpwr.n50 vpwr.n38 4.6505
R517 vpwr.n52 vpwr.n51 4.6505
R518 vpwr.n53 vpwr.n37 4.6505
R519 vpwr.n55 vpwr.n54 4.6505
R520 vpwr.n56 vpwr.n36 4.6505
R521 vpwr.n57 vpwr.n35 4.6505
R522 vpwr.n61 vpwr.n60 4.6505
R523 vpwr.n62 vpwr.n34 4.6505
R524 vpwr.n64 vpwr.n63 4.6505
R525 vpwr.n65 vpwr.n33 4.6505
R526 vpwr.n67 vpwr.n66 4.6505
R527 vpwr.n68 vpwr.n32 4.6505
R528 vpwr.n70 vpwr.n69 4.6505
R529 vpwr.n71 vpwr.n30 4.6505
R530 vpwr.n4 vpwr 4.53383
R531 vpwr.n46 vpwr.n40 4.07323
R532 vpwr.n73 vpwr.n72 3.93272
R533 vpwr.n60 vpwr.n59 3.76521
R534 vpwr.n5 vpwr 3.11401
R535 vpwr.n17 vpwr.n15 3.0725
R536 vpwr.n27 vpwr.n26 2.91783
R537 vpwr.n12 vpwr 2.36657
R538 vpwr.n28 vpwr 1.89029
R539 vpwr.n5 vpwr.n1 1.55726
R540 vpwr.n10 vpwr.n9 1.55726
R541 vpwr.n8 vpwr.n1 1.38428
R542 vpwr.n9 vpwr.n8 1.38428
R543 vpwr.n10 vpwr 1.38428
R544 vpwr.n17 vpwr.n16 1.2805
R545 vpwr.n77 vpwr.n76 0.711611
R546 vpwr.n12 vpwr 0.580857
R547 vpwr.n29 vpwr.n28 0.5255
R548 vpwr.n75 vpwr 0.223
R549 vpwr.n3 vpwr 0.196446
R550 vpwr.n20 vpwr 0.171696
R551 vpwr.n47 vpwr.n42 0.144332
R552 vpwr.n73 vpwr.n30 0.138831
R553 vpwr.n48 vpwr.n47 0.120292
R554 vpwr.n48 vpwr.n38 0.120292
R555 vpwr.n52 vpwr.n38 0.120292
R556 vpwr.n53 vpwr.n52 0.120292
R557 vpwr.n54 vpwr.n53 0.120292
R558 vpwr.n54 vpwr.n36 0.120292
R559 vpwr.n36 vpwr.n35 0.120292
R560 vpwr.n61 vpwr.n35 0.120292
R561 vpwr.n62 vpwr.n61 0.120292
R562 vpwr.n63 vpwr.n62 0.120292
R563 vpwr.n63 vpwr.n33 0.120292
R564 vpwr.n67 vpwr.n33 0.120292
R565 vpwr.n68 vpwr.n67 0.120292
R566 vpwr.n69 vpwr.n68 0.120292
R567 vpwr.n69 vpwr.n30 0.120292
R568 vpwr.n74 vpwr.n73 0.107496
R569 vpwr.n20 vpwr.n19 0.0901739
R570 vpwr vpwr.n83 0.0634013
R571 vpwr.n27 vpwr 0.063
R572 vpwr.n21 vpwr.n20 0.0500874
R573 vpwr.n13 vpwr.n12 0.0466957
R574 vpwr.n24 vpwr.n23 0.0435328
R575 vpwr.n83 vpwr.n29 0.039096
R576 vpwr.n18 vpwr.n13 0.0331087
R577 vpwr.n83 vpwr.n82 0.0287348
R578 vpwr.n3 vpwr.n2 0.02675
R579 vpwr vpwr.n11 0.0255
R580 vpwr.n22 vpwr.n21 0.0213989
R581 vpwr.n78 vpwr.n75 0.0207266
R582 vpwr.n26 vpwr.n25 0.018111
R583 vpwr.n74 vpwr 0.0174271
R584 vpwr vpwr.n74 0.01675
R585 vpwr.n19 vpwr.n18 0.014087
R586 vpwr.n24 vpwr.n22 0.0127951
R587 vpwr.n11 vpwr.n0 0.01175
R588 vpwr.n2 vpwr.n0 0.0105
R589 vpwr.n81 vpwr.n80 0.009875
R590 vpwr vpwr.n3 0.00725676
R591 vpwr.n23 vpwr 0.00459836
R592 vpwr.n79 vpwr.n78 0.00412592
R593 vpwr.n80 vpwr.n79 0.003625
R594 vpwr.n82 vpwr.n81 0.00196888
R595 vpwr.n26 vpwr.n24 0.0016109
R596 vpwr.n78 vpwr.n77 0.00154933
R597 vpwr.n28 vpwr.n27 0.000500433
R598 buffer_0.a.n6 buffer_0.a.t17 377.647
R599 buffer_0.a.n6 buffer_0.a.t16 376.93
R600 buffer_0.a.n13 buffer_0.a.t13 314.055
R601 buffer_0.a.t5 buffer_0.a.n6 42.2586
R602 buffer_0.a.n7 buffer_0.a.t5 40.2461
R603 buffer_0.a.n1 buffer_0.a.t11 39.5847
R604 buffer_0.a.n11 buffer_0.a.t3 39.5292
R605 buffer_0.a.n9 buffer_0.a.t7 39.5292
R606 buffer_0.a.n8 buffer_0.a.t9 39.5292
R607 buffer_0.a.n7 buffer_0.a.t1 39.5292
R608 buffer_0.a.n2 buffer_0.a.t12 28.5655
R609 buffer_0.a.n2 buffer_0.a.t4 28.5655
R610 buffer_0.a.n3 buffer_0.a.t2 28.5655
R611 buffer_0.a.n3 buffer_0.a.t6 28.5655
R612 buffer_0.a.n4 buffer_0.a.t8 28.5655
R613 buffer_0.a.n4 buffer_0.a.t10 28.5655
R614 buffer_0.a.n13 buffer_0.a.t15 13.2078
R615 buffer_0.a.n0 buffer_0.a.t0 13.2005
R616 buffer_0.a.n0 buffer_0.a.t14 13.2005
R617 buffer_0.a.n5 buffer_0.a.n3 1.62643
R618 buffer_0.a.n10 buffer_0.a.n5 1.438
R619 buffer_0.a.n10 buffer_0.a.n9 1.06207
R620 buffer_0.a.n12 buffer_0.a.n11 1.01015
R621 buffer_0.a.n8 buffer_0.a.n7 0.717388
R622 buffer_0.a.n9 buffer_0.a.n8 0.717388
R623 buffer_0.a buffer_0.a.n0 0.677588
R624 buffer_0.a buffer_0.a.n1 0.45343
R625 buffer_0.a.n5 buffer_0.a.n4 0.157684
R626 buffer_0.a.n0 buffer_0.a.n13 0.119008
R627 buffer_0.a.n11 buffer_0.a.n10 0.0949882
R628 buffer_0.a.n1 buffer_0.a.n12 0.0588333
R629 buffer_0.a.n1 buffer_0.a.n2 0.0587685
R630 sensor_0.b.t8 sensor_0.b.t0 74.8549
R631 sensor_0.b.t6 sensor_0.b.t8 74.8549
R632 sensor_0.b.t14 sensor_0.b.t6 74.8549
R633 sensor_0.b.t10 sensor_0.b.t2 74.8549
R634 sensor_0.b.t4 sensor_0.b.t10 74.8549
R635 sensor_0.b.t12 sensor_0.b.t4 74.8549
R636 sensor_0.b.t24 sensor_0.b.t32 74.8549
R637 sensor_0.b.t31 sensor_0.b.t24 74.8549
R638 sensor_0.b.t23 sensor_0.b.t31 74.8549
R639 sensor_0.b.t34 sensor_0.b.t26 74.8549
R640 sensor_0.b.t21 sensor_0.b.t34 74.8549
R641 sensor_0.b.t29 sensor_0.b.t21 74.8549
R642 sensor_0.b.t27 sensor_0.b.t20 74.8549
R643 sensor_0.b.t28 sensor_0.b.t27 74.8549
R644 sensor_0.b.t35 sensor_0.b.t28 74.8549
R645 sensor_0.b.t22 sensor_0.b.t30 74.8549
R646 sensor_0.b.t33 sensor_0.b.t22 74.8549
R647 sensor_0.b.t25 sensor_0.b.t33 74.8549
R648 sensor_0.b.n7 sensor_0.b.t25 38.3763
R649 sensor_0.b.n11 sensor_0.b.t14 37.3627
R650 sensor_0.b.n10 sensor_0.b.t12 37.3602
R651 sensor_0.b.n9 sensor_0.b.t23 37.3602
R652 sensor_0.b.n8 sensor_0.b.t29 37.3602
R653 sensor_0.b.n7 sensor_0.b.t35 37.3602
R654 sensor_0.b.n12 sensor_0.b.t1 18.2715
R655 sensor_0.b.n3 sensor_0.b.t3 18.1717
R656 sensor_0.b.n14 sensor_0.b.t15 17.427
R657 sensor_0.b.n13 sensor_0.b.t7 17.4116
R658 sensor_0.b.n3 sensor_0.b.t11 17.4101
R659 sensor_0.b.n12 sensor_0.b.t9 17.4101
R660 sensor_0.b.n4 sensor_0.b.t5 17.4058
R661 sensor_0.b.n5 sensor_0.b.t13 17.4056
R662 sensor_0.b.n0 sensor_0.b.t19 14.283
R663 sensor_0.b.n0 sensor_0.b.t18 14.283
R664 sensor_0.b.n1 sensor_0.b.t16 14.283
R665 sensor_0.b.n1 sensor_0.b.t17 14.283
R666 sensor_0.b.n6 sensor_0.b.n5 3.22928
R667 sensor_0.b.n6 sensor_0.b.n2 2.2255
R668 sensor_0.b.n11 sensor_0.b.n10 1.01759
R669 sensor_0.b.n8 sensor_0.b.n7 1.01657
R670 sensor_0.b.n9 sensor_0.b.n8 1.01657
R671 sensor_0.b.n10 sensor_0.b.n9 1.01657
R672 sensor_0.b.n13 sensor_0.b.n12 0.865287
R673 sensor_0.b sensor_0.b.n15 0.851048
R674 sensor_0.b.n14 sensor_0.b.n13 0.777059
R675 sensor_0.b.n5 sensor_0.b.n4 0.718555
R676 sensor_0.b.n4 sensor_0.b.n3 0.710921
R677 sensor_0.b.n2 sensor_0.b.n0 0.49917
R678 sensor_0.b sensor_0.b.n6 0.341125
R679 sensor_0.b.n15 sensor_0.b.n14 0.325292
R680 sensor_0.b.n15 sensor_0.b.n11 0.202053
R681 sensor_0.b.n2 sensor_0.b.n1 0.17167
R682 sensor_0.a.n2 sensor_0.a.t15 64.1667
R683 sensor_0.a.n0 sensor_0.a.t2 63.6292
R684 sensor_0.a.n4 sensor_0.a.t13 63.6292
R685 sensor_0.a.n3 sensor_0.a.t12 63.6292
R686 sensor_0.a.n2 sensor_0.a.t14 63.6292
R687 sensor_0.a.n1 sensor_0.a.t0 63.6275
R688 sensor_0.a.n8 sensor_0.a.t6 18.2715
R689 sensor_0.a.n5 sensor_0.a.t11 18.2714
R690 sensor_0.a.n10 sensor_0.a.t9 17.4132
R691 sensor_0.a.n7 sensor_0.a.t4 17.4132
R692 sensor_0.a.n6 sensor_0.a.t7 17.4116
R693 sensor_0.a.n8 sensor_0.a.t10 17.4101
R694 sensor_0.a.n5 sensor_0.a.t8 17.4101
R695 sensor_0.a.n9 sensor_0.a.t5 17.4057
R696 sensor_0.a.n1 sensor_0.a.t1 14.5343
R697 sensor_0.a.n0 sensor_0.a.t3 14.2976
R698 sensor_0.a sensor_0.a.n11 1.63801
R699 sensor_0.a.n11 sensor_0.a.n7 1.541
R700 sensor_0.a.n11 sensor_0.a.n10 1.541
R701 sensor_0.a.n10 sensor_0.a.n9 0.873387
R702 sensor_0.a.n6 sensor_0.a.n5 0.865287
R703 sensor_0.a.n7 sensor_0.a.n6 0.864262
R704 sensor_0.a.n9 sensor_0.a.n8 0.848309
R705 sensor_0.a.n3 sensor_0.a.n2 0.538
R706 sensor_0.a.n4 sensor_0.a.n3 0.538
R707 sensor_0.a.n0 sensor_0.a.n4 0.488
R708 sensor_0.a.n1 sensor_0.a.n0 0.29354
R709 sensor_0.a sensor_0.a.n1 0.28675
R710 buffer_0.b.n6 buffer_0.b.t17 377.466
R711 buffer_0.b.n6 buffer_0.b.t16 376.93
R712 buffer_0.b.n16 buffer_0.b.t0 313.991
R713 buffer_0.b.t7 buffer_0.b.n6 41.3792
R714 buffer_0.b.n7 buffer_0.b.t7 40.2104
R715 buffer_0.b.n11 buffer_0.b.t4 28.6605
R716 buffer_0.b.n0 buffer_0.b.t10 28.5655
R717 buffer_0.b.n0 buffer_0.b.t3 28.5655
R718 buffer_0.b.n2 buffer_0.b.t8 28.5655
R719 buffer_0.b.n2 buffer_0.b.t12 28.5655
R720 buffer_0.b.n3 buffer_0.b.t6 28.5655
R721 buffer_0.b.n3 buffer_0.b.t14 28.5655
R722 buffer_0.b.n11 buffer_0.b.t2 26.2653
R723 buffer_0.b.n10 buffer_0.b.t9 26.2652
R724 buffer_0.b.n9 buffer_0.b.t13 26.2652
R725 buffer_0.b.n8 buffer_0.b.t5 26.2652
R726 buffer_0.b.n7 buffer_0.b.t11 26.2652
R727 buffer_0.b.n15 buffer_0.b.t15 13.2053
R728 buffer_0.b.n15 buffer_0.b.t1 6.63265
R729 buffer_0.b.n4 buffer_0.b.n2 1.62544
R730 buffer_0.b.n5 buffer_0.b.n4 1.44539
R731 buffer_0.b.n1 buffer_0.b.n10 0.825504
R732 buffer_0.b.n8 buffer_0.b.n7 0.718158
R733 buffer_0.b.n9 buffer_0.b.n8 0.718158
R734 buffer_0.b.n10 buffer_0.b.n9 0.718158
R735 buffer_0.b buffer_0.b.n16 0.594255
R736 buffer_0.b buffer_0.b.n14 0.562809
R737 buffer_0.b.n13 buffer_0.b.n12 0.188
R738 buffer_0.b.n4 buffer_0.b.n3 0.156686
R739 buffer_0.b.n12 buffer_0.b.n1 0.10675
R740 buffer_0.b.n13 buffer_0.b.n5 0.104667
R741 buffer_0.b.n16 buffer_0.b.n15 0.0678366
R742 buffer_0.b.n14 buffer_0.b.n0 0.0624088
R743 buffer_0.b.n1 buffer_0.b.n11 0.0623624
R744 buffer_0.b.n0 buffer_0.b.n13 0.0505
R745 out_buff.n4 out_buff.t7 377.192
R746 out_buff.n1 out_buff.t5 377.175
R747 out_buff.n6 out_buff.t11 317.7
R748 out_buff.n13 out_buff.t4 9.50808
R749 out_buff.n12 out_buff 6.13573
R750 out_buff.n9 out_buff.t9 5.53268
R751 out_buff.n7 out_buff.t3 3.4805
R752 out_buff.n7 out_buff.t2 3.4805
R753 out_buff.n12 out_buff.n11 2.388
R754 out_buff.n5 out_buff.n4 2.02858
R755 out_buff.n2 out_buff.n1 2.00736
R756 out_buff.n3 out_buff.t1 1.90483
R757 out_buff.n3 out_buff.t8 1.90483
R758 out_buff.n0 out_buff.t6 1.90483
R759 out_buff.n0 out_buff.t0 1.90483
R760 out_buff.n6 out_buff.t10 1.78624
R761 out_buff.n8 out_buff.n7 1.58206
R762 out_buff.n13 out_buff.n12 1.11925
R763 out_buff.n10 out_buff.n9 0.80675
R764 out_buff.n9 out_buff.n8 0.770812
R765 out_buff.n11 out_buff.n10 0.722063
R766 out_buff.n10 out_buff.n2 0.182565
R767 out_buff.n9 out_buff.n5 0.182565
R768 out_buff.n11 out_buff 0.06175
R769 out_buff out_buff.n13 0.05675
R770 out_buff.n5 out_buff.n3 0.00195207
R771 out_buff.n2 out_buff.n0 0.00195207
R772 out_buff.n8 out_buff.n6 0.000558569
R773 vd.n61 vd.n43 11483
R774 vd.n56 vd.n43 11371.8
R775 vd.n64 vd.n42 10557.3
R776 vd.n53 vd.n52 10507.9
R777 vd.n45 vd.n42 8128.24
R778 vd.n52 vd.n47 8092.94
R779 vd.n56 vd.n47 6967.06
R780 vd.n61 vd.n45 6931.77
R781 vd.n64 vd.n40 6349.41
R782 vd.n53 vd.n40 6345.88
R783 vd.n18 vd.n15 2142.35
R784 vd.n60 vd.n58 1224.85
R785 vd.n58 vd.n57 1212.99
R786 vd.n22 vd.n16 1164.71
R787 vd.n24 vd.n12 1164.71
R788 vd.n65 vd.n41 1126.12
R789 vd.n50 vd.n39 1120.84
R790 vd.n24 vd.n13 977.648
R791 vd.n22 vd.n15 952.942
R792 vd.n59 vd.n41 867.013
R793 vd.n50 vd.n46 863.247
R794 vd.n57 vd.n46 743.154
R795 vd.n60 vd.n59 739.389
R796 vd.n66 vd.n65 647.907
R797 vd.n66 vd.n39 647.529
R798 vd.t63 vd.t6 331.216
R799 vd.t6 vd.t12 331.216
R800 vd.t12 vd.t10 331.216
R801 vd.t10 vd.t1 331.216
R802 vd.t1 vd.t8 331.216
R803 vd.t8 vd.t5 331.216
R804 vd.t41 vd.t39 331.216
R805 vd.t39 vd.t42 331.216
R806 vd.t42 vd.t33 331.216
R807 vd.t33 vd.t31 331.216
R808 vd.t31 vd.t29 331.216
R809 vd.t29 vd.t66 331.216
R810 vd.n20 vd.n19 228.518
R811 vd.n19 vd.n10 228.518
R812 vd.n48 vd.t41 228.514
R813 vd.t5 vd.n49 210.542
R814 vd.n137 vd.n134 206.306
R815 vd.n105 vd.n104 168.66
R816 vd.t55 vd.n118 156.245
R817 vd.n23 vd.t16 144.606
R818 vd.n100 vd.t49 143.697
R819 vd.n122 vd.t23 143.697
R820 vd.n144 vd.n141 142.306
R821 vd.n18 vd.n17 135.465
R822 vd.n124 vd.n121 126.871
R823 vd.n97 vd.n96 111.421
R824 vd.n25 vd.n10 104.282
R825 vd.n21 vd.n20 101.647
R826 vd.n142 vd.t46 86.6752
R827 vd.n105 vd.n99 85.0829
R828 vd.n135 vd.t59 71.8492
R829 vd.t37 vd.t0 70.1694
R830 vd.t35 vd.t52 70.1694
R831 vd.t27 vd.t3 70.0291
R832 vd.t14 vd.t28 70.0291
R833 vd.n62 vd.t0 68.5376
R834 vd.n100 vd.t70 65.0065
R835 vd.n107 vd.t58 63.9214
R836 vd.n93 vd.t69 63.8352
R837 vd.t52 vd.n42 63.6434
R838 vd.n113 vd.t54 63.6292
R839 vd.n55 vd.t28 63.5148
R840 vd.n137 vd.n131 63.2476
R841 vd.n52 vd.t27 62.9732
R842 vd.n142 vd.t47 60.4447
R843 vd.t46 vd.t50 58.1638
R844 vd.t59 vd.t22 58.1638
R845 vd.n129 vd.t44 42.1974
R846 vd.n132 vd.t21 42.1974
R847 vd.n81 vd.t62 39.5312
R848 vd.n71 vd.t65 39.5292
R849 vd.n49 vd.n48 38.514
R850 vd.n44 vd.t35 37.5327
R851 vd.t3 vd.n51 35.2862
R852 vd.n51 vd.t14 34.7434
R853 vd.n44 vd.t37 32.6372
R854 vd.n26 vd.n25 31.105
R855 vd.t64 vd.n81 28.7267
R856 vd.n71 vd.t68 28.6459
R857 vd.n86 vd.t2 28.5655
R858 vd.n86 vd.t9 28.5655
R859 vd.n82 vd.t64 28.5655
R860 vd.n82 vd.t7 28.5655
R861 vd.n84 vd.t13 28.5655
R862 vd.n84 vd.t11 28.5655
R863 vd.n68 vd.t40 28.5655
R864 vd.n68 vd.t43 28.5655
R865 vd.n70 vd.t30 28.5655
R866 vd.n70 vd.t67 28.5655
R867 vd.n73 vd.t34 28.5655
R868 vd.n73 vd.t32 28.5655
R869 vd.n102 vd.t48 28.5119
R870 vd.n21 vd.n4 27.9188
R871 vd.n115 vd.n110 24.5501
R872 vd.n26 vd.n9 22.401
R873 vd.n34 vd.n33 22.4005
R874 vd.n9 vd.n7 22.4005
R875 vd.n55 vd.n54 21.216
R876 vd.n119 vd.t55 21.0989
R877 vd.t44 vd.t19 19.3883
R878 vd.n35 vd.n4 19.201
R879 vd.n35 vd.n34 19.2005
R880 vd.n135 vd.t20 17.1073
R881 vd.n54 vd.n53 16.7426
R882 vd.n63 vd.t66 16.3842
R883 vd.n63 vd.n62 16.211
R884 vd.n106 vd.t45 14.575
R885 vd.n92 vd.t51 14.5025
R886 vd.n112 vd.t56 14.4041
R887 vd.n94 vd.t71 14.2873
R888 vd.n92 vd.t72 14.2873
R889 vd.n108 vd.t61 14.2873
R890 vd.n106 vd.t60 14.2873
R891 vd.n110 vd.t57 14.2867
R892 vd.n111 vd.t24 14.283
R893 vd.n111 vd.t26 14.283
R894 vd.n54 vd.t63 12.5482
R895 vd.t70 vd.t18 11.4051
R896 vd.n11 vd.n7 10.5605
R897 vd.n33 vd.n6 9.6005
R898 vd.n2 vd.t53 9.5742
R899 vd.n30 vd.t17 9.52337
R900 vd.n115 vd.n114 9.3005
R901 vd.n64 vd.n63 7.64222
R902 vd.n116 vd.n115 4.5005
R903 vd.n75 vd.n67 4.5005
R904 vd vd.n38 4.16717
R905 vd.n149 vd.n148 3.79434
R906 vd.n88 vd.n80 3.54402
R907 vd.n79 vd.n78 3.47391
R908 vd.n122 vd.t25 3.42187
R909 vd.n11 vd.n6 2.2405
R910 vd.n80 vd.t4 1.90483
R911 vd.n80 vd.t15 1.90483
R912 vd.n78 vd.t38 1.90483
R913 vd.n78 vd.t36 1.90483
R914 vd vd.n116 1.83279
R915 vd.n91 vd 1.73266
R916 vd.n85 vd.n83 1.56925
R917 vd.n74 vd.n72 1.5417
R918 vd.n87 vd.n85 1.44593
R919 vd.n75 vd.n74 1.38331
R920 vd.n147 vd.n94 0.881455
R921 vd.n148 vd.n147 0.834744
R922 vd.n112 vd.n111 0.721906
R923 vd.n83 vd.n81 0.686006
R924 vd.n113 vd.n112 0.608294
R925 vd.n126 vd.n108 0.59946
R926 vd.n146 vd.n145 0.5755
R927 vd.n89 vd.n79 0.497524
R928 vd.n145 vd.n138 0.488
R929 vd.n126 vd.n125 0.463
R930 vd.n89 vd.n88 0.4255
R931 vd.n88 vd.n87 0.424134
R932 vd.n148 vd.n91 0.328325
R933 vd.n79 vd.n77 0.313286
R934 vd.n125 vd 0.2755
R935 vd.n138 vd.n126 0.238
R936 vd.n150 vd.n149 0.2005
R937 vd.n85 vd.n84 0.157684
R938 vd.n74 vd.n73 0.156686
R939 vd.n28 vd.n27 0.146341
R940 vd.n28 vd.n3 0.146333
R941 vd.n107 vd.n106 0.134875
R942 vd.n108 vd.n107 0.134875
R943 vd.n22 vd.n21 0.130052
R944 vd.n23 vd.n22 0.130052
R945 vd.n38 vd.n3 0.1255
R946 vd.n150 vd 0.1255
R947 vd.n110 vd.n109 0.122252
R948 vd.n114 vd.n113 0.116172
R949 vd.n94 vd.n93 0.115679
R950 vd.n93 vd.n92 0.115679
R951 vd.n25 vd.n24 0.107375
R952 vd.n24 vd.n23 0.107375
R953 vd.n91 vd 0.100725
R954 vd.n150 vd.n2 0.0822638
R955 vd.n72 vd.n71 0.0791768
R956 vd.n0 vd.t73 0.0686501
R957 vd.n1 vd.n0 0.06865
R958 vd.n72 vd.n70 0.0493677
R959 vd.n76 vd.n75 0.0489375
R960 vd.n83 vd.n82 0.0461626
R961 vd.n32 vd.n5 0.0456031
R962 vd.n29 vd.n8 0.0456031
R963 vd.n27 vd.n8 0.0456031
R964 vd.n37 vd.n36 0.0391598
R965 vd.n36 vd.n5 0.0391598
R966 vd.n149 vd 0.0372647
R967 vd.n20 vd.n15 0.0349892
R968 vd.n15 vd.t16 0.0349892
R969 vd.n13 vd.n10 0.0349892
R970 vd vd.n90 0.0347717
R971 vd.n17 vd.n13 0.0333079
R972 vd.n99 vd.n98 0.0307238
R973 vd.n98 vd.n97 0.0302348
R974 vd.n30 vd.n29 0.0217629
R975 vd.n69 vd.n68 0.0200317
R976 vd.n32 vd.n31 0.0198299
R977 vd.n77 vd.n67 0.01975
R978 vd.n116 vd.n109 0.0176875
R979 vd.n121 vd.n120 0.0175052
R980 vd.n120 vd.n119 0.0175052
R981 vd.n141 vd.n140 0.0150968
R982 vd.n140 vd.n139 0.0150968
R983 vd.n87 vd.n86 0.0148061
R984 vd.n69 vd.n67 0.0141783
R985 vd vd.n150 0.013
R986 vd.n14 vd.n12 0.0125538
R987 vd.n104 vd.n103 0.0122827
R988 vd.n103 vd.n102 0.0122827
R989 vd.n12 vd.n11 0.0120596
R990 vd.n114 vd.n109 0.009875
R991 vd.n134 vd.n133 0.00973799
R992 vd.n133 vd.n132 0.00973799
R993 vd.n2 vd.n1 0.00846782
R994 vd.n76 vd.n69 0.0083125
R995 vd.n147 vd.n146 0.00675
R996 vd.n19 vd.n18 0.00627981
R997 vd.n31 vd.n30 0.00501031
R998 vd.n47 vd.n46 0.00431884
R999 vd.n51 vd.n47 0.00431884
R1000 vd.n59 vd.n45 0.00425193
R1001 vd.n45 vd.n44 0.00425193
R1002 vd.n144 vd.n143 0.00391284
R1003 vd.n143 vd.n142 0.00391284
R1004 vd.n137 vd.n136 0.00391284
R1005 vd.n136 vd.n135 0.00391284
R1006 vd.n124 vd.n123 0.00391284
R1007 vd.n123 vd.n122 0.00391284
R1008 vd.n105 vd.n101 0.00391284
R1009 vd.n101 vd.n100 0.00391284
R1010 vd.n65 vd.n64 0.00389051
R1011 vd.n53 vd.n39 0.00389051
R1012 vd.n118 vd.n117 0.00347027
R1013 vd.n96 vd.n95 0.00347027
R1014 vd.n17 vd.t16 0.00318081
R1015 vd.n131 vd.n130 0.00275116
R1016 vd.n130 vd.n129 0.00275116
R1017 vd.n61 vd.n60 0.0021559
R1018 vd.n62 vd.n61 0.0021559
R1019 vd.n57 vd.n56 0.00213065
R1020 vd.n56 vd.n55 0.00213065
R1021 vd.n90 vd.n66 0.00200289
R1022 vd.n16 vd.n14 0.0018171
R1023 vd.n42 vd.n41 0.00181202
R1024 vd.n52 vd.n50 0.00181202
R1025 vd.n58 vd.n43 0.0017783
R1026 vd.n49 vd.n43 0.0017783
R1027 vd.n129 vd.n128 0.00162558
R1028 vd.n128 vd.n127 0.00162558
R1029 vd.n16 vd.n6 0.00131751
R1030 vd.n31 vd.n6 0.00131744
R1031 vd.n36 vd.n35 0.00119114
R1032 vd.n37 vd.n4 0.00101609
R1033 vd.n77 vd.n76 0.00100557
R1034 vd.n90 vd.n89 0.00100109
R1035 vd.n23 vd.n14 0.00100038
R1036 vd.n27 vd.n26 0.00100009
R1037 vd.n66 vd.n40 0.000827345
R1038 vd.n48 vd.n40 0.000827345
R1039 vd.n9 vd.n8 0.000659706
R1040 vd.n33 vd.n32 0.000659706
R1041 vd.n34 vd.n5 0.000543686
R1042 vd.n29 vd.n7 0.000543686
R1043 vd.n145 vd.n144 0.000532663
R1044 vd.n138 vd.n137 0.000532663
R1045 vd.n125 vd.n124 0.000532663
R1046 vd.n146 vd.n105 0.000532663
R1047 vd.n38 vd.n37 0.000507883
R1048 vd.n5 vd.n3 0.000507883
R1049 vd.n29 vd.n28 0.000507883
R1050 vd.n0 vd.t75 0.000500086
R1051 vd.n1 vd.t74 0.000500086
R1052 vtd.n7 vtd.t29 64.6821
R1053 vtd.n8 vtd.t27 64.3461
R1054 vtd.n4 vtd.t24 63.6317
R1055 vtd.n9 vtd.t26 63.6292
R1056 vtd.n8 vtd.t28 63.6292
R1057 vtd.n17 vtd.t2 63.6292
R1058 vtd.n2 vtd.t10 63.6292
R1059 vtd.n18 vtd.t14 63.6292
R1060 vtd.n1 vtd.t8 63.6292
R1061 vtd.n19 vtd.t0 63.6292
R1062 vtd.n0 vtd.t6 63.6292
R1063 vtd.n6 vtd.t12 63.6292
R1064 vtd.n3 vtd.t4 63.6275
R1065 vtd.n13 vtd.t20 18.2948
R1066 vtd.n10 vtd.t17 18.1899
R1067 vtd.n10 vtd.t21 17.4187
R1068 vtd.n13 vtd.t16 17.4177
R1069 vtd.n11 vtd.t18 17.4156
R1070 vtd.n14 vtd.t23 17.4136
R1071 vtd.n12 vtd.t22 17.4125
R1072 vtd.n15 vtd.t19 17.4115
R1073 vtd.n3 vtd.t5 14.3559
R1074 vtd.n17 vtd.t3 14.3555
R1075 vtd.n2 vtd.t15 14.283
R1076 vtd.n2 vtd.t11 14.283
R1077 vtd.n1 vtd.t1 14.283
R1078 vtd.n1 vtd.t9 14.283
R1079 vtd.n0 vtd.t13 14.283
R1080 vtd.n0 vtd.t7 14.283
R1081 vtd.n7 vtd.t25 13.7801
R1082 vtd.n16 vtd.n15 2.14635
R1083 vtd.n3 vtd.n16 1.54335
R1084 vtd vtd.n20 1.22372
R1085 vtd.n16 vtd.n12 1.09526
R1086 vtd.n20 vtd.n3 0.981002
R1087 vtd.n15 vtd.n14 0.8755
R1088 vtd.n14 vtd.n13 0.8755
R1089 vtd.n5 vtd.n7 0.832184
R1090 vtd.n11 vtd.n10 0.769433
R1091 vtd.n12 vtd.n11 0.769356
R1092 vtd.n9 vtd.n8 0.717388
R1093 vtd.n4 vtd.n9 0.708453
R1094 vtd.n20 vtd.n5 0.438348
R1095 vtd.n3 vtd.n6 0.140567
R1096 vtd.n18 vtd.n2 0.140142
R1097 vtd.n19 vtd.n1 0.140142
R1098 vtd.n6 vtd.n0 0.140142
R1099 vtd.n0 vtd.n19 0.134875
R1100 vtd.n1 vtd.n18 0.134875
R1101 vtd.n2 vtd.n17 0.134875
R1102 vtd.n5 vtd.n4 0.114328
R1103 buffer_0.d.n9 buffer_0.d.t2 377.216
R1104 buffer_0.d.n8 buffer_0.d.t0 377.163
R1105 buffer_0.d.n2 buffer_0.d.t12 134.298
R1106 buffer_0.d.n4 buffer_0.d.t5 133.787
R1107 buffer_0.d.n3 buffer_0.d.t7 133.761
R1108 buffer_0.d.n2 buffer_0.d.t13 133.761
R1109 buffer_0.d.n1 buffer_0.d.t4 5.55126
R1110 buffer_0.d.n6 buffer_0.d.t8 3.4805
R1111 buffer_0.d.n6 buffer_0.d.t6 3.4805
R1112 buffer_0.d buffer_0.d.n7 3.10062
R1113 buffer_0.d.n1 buffer_0.d.n9 2.02586
R1114 buffer_0.d.n0 buffer_0.d.n8 1.99422
R1115 buffer_0.d.n5 buffer_0.d.t9 1.91167
R1116 buffer_0.d.n0 buffer_0.d.t11 1.9057
R1117 buffer_0.d.n1 buffer_0.d.t10 1.90483
R1118 buffer_0.d.n1 buffer_0.d.t3 1.90483
R1119 buffer_0.d.n0 buffer_0.d.t1 1.42659
R1120 buffer_0.d buffer_0.d.n0 0.77675
R1121 buffer_0.d.n0 buffer_0.d.n1 0.648539
R1122 buffer_0.d.n3 buffer_0.d.n2 0.538
R1123 buffer_0.d.n4 buffer_0.d.n3 0.394346
R1124 buffer_0.d.n7 buffer_0.d.n6 0.151643
R1125 buffer_0.d.n5 buffer_0.d.n4 0.0558728
R1126 buffer_0.d.n7 buffer_0.d.n5 0.0333947
R1127 ib.n0 ib.t5 38.0465
R1128 ib.n0 ib.t0 37.3602
R1129 ib.n4 ib.t2 18.7496
R1130 ib.n4 ib.t4 17.4934
R1131 ib.n1 ib.t1 17.4005
R1132 ib.n1 ib.t3 17.4005
R1133 ib.n9 ib.n8 5.70556
R1134 ib.n3 ib.n2 1.98477
R1135 ib.n8 ib.n0 0.247263
R1136 ib.n10 ib 0.129406
R1137 ib.n9 ib 0.1205
R1138 ib.n5 ib.n4 0.102062
R1139 ib ib.n10 0.0605
R1140 ib.n8 ib.n7 0.059593
R1141 ib.n7 ib.n6 0.0239375
R1142 ib.n6 ib.n3 0.0166802
R1143 ib.n6 ib.n5 0.003625
R1144 ib.n3 ib.n1 0.00322924
R1145 ib.n10 ib.n9 0.00114405
R1146 vts.n23 vts.n18 761.601
R1147 vts.n24 vts.n23 641.883
R1148 vts.t18 vts.t4 333.303
R1149 vts.n35 vts.t25 325.759
R1150 vts.n17 vts.t22 262.014
R1151 vts.n26 vts.t18 237.054
R1152 vts.t4 vts.t2 229.925
R1153 vts.t15 vts.t0 229.925
R1154 vts.t13 vts.t11 229.925
R1155 vts.t11 vts.t9 229.925
R1156 vts.t9 vts.t7 229.925
R1157 vts.n21 vts.t15 130.113
R1158 vts.n21 vts.t13 99.8129
R1159 vts.n11 vts.t17 63.6292
R1160 vts.n4 vts.t21 63.6292
R1161 vts.n31 vts.t6 16.8006
R1162 vts.n5 vts.t23 14.4639
R1163 vts.n10 vts.t20 14.4362
R1164 vts.n12 vts.t19 14.4313
R1165 vts.n4 vts.t24 14.3697
R1166 vts.n0 vts.t5 14.283
R1167 vts.n0 vts.t3 14.283
R1168 vts.n1 vts.t1 14.283
R1169 vts.n1 vts.t16 14.283
R1170 vts.n2 vts.t14 14.283
R1171 vts.n2 vts.t12 14.283
R1172 vts.n3 vts.t10 14.283
R1173 vts.n3 vts.t8 14.283
R1174 vts.n36 vts 3.48645
R1175 vts.n36 vts.n35 1.21925
R1176 vts vts.n34 0.8255
R1177 vts.n9 vts.n8 0.6455
R1178 vts.n8 vts.n7 0.6455
R1179 vts.n7 vts.n6 0.6455
R1180 vts.n6 vts.n5 0.450361
R1181 vts.n10 vts.n9 0.440551
R1182 vts vts.n36 0.26925
R1183 vts.n30 vts.n12 0.0947919
R1184 vts.n5 vts.n4 0.0741592
R1185 vts.n11 vts.n10 0.0682354
R1186 vts.n12 vts.n11 0.0634447
R1187 vts.n35 vts 0.058
R1188 vts.n34 vts.n33 0.05093
R1189 vts.n25 vts.n24 0.0426316
R1190 vts.n26 vts.n25 0.0426316
R1191 vts.n16 vts.n15 0.0175052
R1192 vts.n26 vts.n16 0.0175052
R1193 vts.n9 vts.n0 0.0129196
R1194 vts.n8 vts.n1 0.0129196
R1195 vts.n7 vts.n2 0.0129196
R1196 vts.n6 vts.n3 0.0129196
R1197 vts.n27 vts.n14 0.011183
R1198 vts.n14 vts.n13 0.0106833
R1199 vts.n28 vts.n27 0.0075124
R1200 vts.n29 vts.n28 0.00701261
R1201 vts.n18 vts.n17 0.00559165
R1202 vts.n23 vts.n22 0.00192573
R1203 vts.n22 vts.n21 0.00192573
R1204 vts.n20 vts.n19 0.00192573
R1205 vts.n21 vts.n20 0.00192573
R1206 vts.n33 vts.n32 0.00151802
R1207 vts.n32 vts.n30 0.00150795
R1208 vts.n27 vts.n26 0.00100013
R1209 vts.n30 vts.n29 0.00100001
R1210 vts.n32 vts.n31 0.001
R1211 clk.n0 clk.t1 294.557
R1212 clk.n0 clk.t0 211.01
R1213 clk.n2 clk.n0 8.28655
R1214 clk.n3 clk 7.73487
R1215 clk.n3 clk.n2 1.82961
R1216 clk.n1 clk 0.981259
R1217 clk.n2 clk.n1 0.848973
R1218 clk clk.n5 0.385917
R1219 clk.n5 clk.n4 0.03175
R1220 clk.n4 clk.n3 0.00111796
R1221 out.n2 out.t0 8.97158
R1222 out.n2 out.n1 2.56714
R1223 out.n0 out.t2 0.506271
R1224 out.n1 out.n0 0.504061
R1225 out out.n2 0.240344
R1226 out.n0 out.t1 0.0277714
R1227 out.n1 out.t3 0.00303875
R1228 out_sigma.n2 out_sigma.t2 394.808
R1229 out_sigma.n0 out_sigma.t1 250.941
R1230 out_sigma out_sigma.t0 144.601
R1231 out_sigma out_sigma.n2 9.0826
R1232 out_sigma.n1 out_sigma.n0 4.66
R1233 out_sigma.n3 out_sigma 4.17039
R1234 out_sigma.n0 out_sigma 3.35288
R1235 out_sigma.n3 out_sigma 3.1826
R1236 out_sigma.n2 out_sigma 0.727062
R1237 out_sigma.n1 out_sigma 0.6255
R1238 out_sigma out_sigma.n3 0.13175
R1239 out_sigma out_sigma.n1 0.063
C0 out_buff a_14882_5320# 0.0014f
C1 a_15546_5320# a_15214_5320# 0.296f
C2 vpwr a_15249_1221# 0.156f
C3 a_16688_5320# sigma-delta_0.x1.Q 0.0032f
C4 clk a_14791_855# 0.00241f
C5 sigma-delta_0.in_int a_15098_3152# 0.0613f
C6 clk a_14600_2320# 1.96e-19
C7 a_15214_5320# sigma-delta_0.in_int 0.00277f
C8 a_16854_3988# a_17020_5320# 0.00434f
C9 clk a_15237_855# 5.33e-20
C10 buffer_0.b buffer_0.a 0.239f
C11 a_14625_855# a_14791_855# 0.906f
C12 a_16445_855# a_14791_855# 2.01e-19
C13 sensor_0.a sensor_0.b 0.821f
C14 buffer_0.b buffer_0.d 0.0351f
C15 a_14625_855# a_14600_2320# 1.68e-19
C16 a_17020_5320# sigma-delta_0.in_int 0.00986f
C17 a_15881_829# vpwr 0.688f
C18 vd a_15214_5320# 0.0598f
C19 a_14625_855# a_15237_855# 0.00134f
C20 out out_sigma 5.44f
C21 out_sigma sigma-delta_0.in_comp 0.0553f
C22 a_15359_1097# a_15706_855# 0.0512f
C23 out_buff a_15380_3988# 5.35e-19
C24 a_14766_3152# a_14932_2320# 0.00938f
C25 a_14600_2320# sigma-delta_0.in_int 0.0164f
C26 a_15430_3152# a_15380_3988# 0.00472f
C27 buffer_0.d buffer_0.a 1.27f
C28 vts sensor_0.d 0.248f
C29 a_15046_855# sigma-delta_0.x1.Q 7.58e-20
C30 a_15815_855# a_14791_855# 2.36e-20
C31 sensor_0.a sensor_0.c 0.997f
C32 sigma-delta_0.x1.D a_15706_855# 9.45e-19
C33 a_15141_855# a_14791_855# 0.23f
C34 vd a_17020_5320# 0.201f
C35 vd a_14791_855# 1.08e-19
C36 a_14550_5320# sigma-delta_0.in_int 0.00283f
C37 a_15141_855# a_15237_855# 0.0138f
C38 a_15098_3152# a_14932_2320# 0.00938f
C39 out a_14882_5320# 0.0019f
C40 sensor_0.c sensor_0.b 0.55f
C41 a_16060_855# sigma-delta_0.x1.Q 6.05e-19
C42 vts ib 1.08f
C43 a_14625_855# a_15596_2320# 1.47e-19
C44 vd a_14550_5320# 0.067f
C45 a_15868_1221# sigma-delta_0.x1.Q 4.53e-20
C46 vd sensor_0.d 0.282f
C47 a_16522_3988# a_16854_3988# 0.303f
C48 out_sigma a_15881_829# 0.00735f
C49 a_15596_2320# sigma-delta_0.in_int 0.00497f
C50 a_14791_855# a_14932_2320# 1.47e-19
C51 a_16688_5320# a_17020_5320# 0.299f
C52 a_14600_2320# a_14932_2320# 0.296f
C53 a_16522_3988# sigma-delta_0.in_int 0.0509f
C54 sigma-delta_0.x1.Q a_15098_3152# 1.13e-19
C55 sigma-delta_0.in_int a_14716_3988# 0.0408f
C56 out_sigma vpwr 1.81f
C57 sigma-delta_0.in_comp a_15706_855# 5.26e-20
C58 a_15141_855# a_15596_2320# 1.87e-19
C59 vd a_15596_2320# 1.16e-19
C60 vd ib 0.0124f
C61 out_buff clk 0.683f
C62 clk a_15359_1097# 1.78e-19
C63 a_15403_855# a_15359_1097# 3.69e-19
C64 vd a_16522_3988# 0.00558f
C65 sigma-delta_0.x1.Q a_17020_5320# 0.00839f
C66 vd a_14716_3988# 0.0021f
C67 a_14791_855# sigma-delta_0.x1.Q 0.00137f
C68 out_buff vts 0.103f
C69 out_buff a_15546_5320# 2.84e-19
C70 clk sigma-delta_0.x1.D 0.00993f
C71 a_15264_2320# sigma-delta_0.in_int 0.00497f
C72 out_buff a_14625_855# 4.76e-19
C73 a_15403_855# sigma-delta_0.x1.D 5.41e-20
C74 a_14625_855# a_15359_1097# 0.0701f
C75 a_15237_855# sigma-delta_0.x1.Q 1.45e-19
C76 sensor_0.d sensor_0.a 0.588f
C77 out_buff a_16024_5320# 3.49e-20
C78 a_14791_855# a_15046_855# 0.0642f
C79 out_buff sigma-delta_0.in_int 0.0662f
C80 a_16356_5320# a_16522_3988# 0.00509f
C81 a_15430_3152# sigma-delta_0.in_int 0.0597f
C82 a_14766_3152# a_15098_3152# 0.296f
C83 a_14625_855# sigma-delta_0.x1.D 0.195f
C84 a_16445_855# sigma-delta_0.x1.D 0.00209f
C85 a_15046_855# a_15237_855# 4.61e-19
C86 a_15881_829# a_15706_855# 0.251f
C87 sigma-delta_0.x1.D sigma-delta_0.in_int 0.0121f
C88 a_14882_5320# a_15048_3988# 0.00482f
C89 a_16522_3988# a_16688_5320# 0.00482f
C90 sensor_0.d sensor_0.b 0.0152f
C91 a_15815_855# a_15359_1097# 4.2e-19
C92 out_buff vd 5.19f
C93 a_15141_855# a_15359_1097# 0.21f
C94 vd a_6126_29386# 0.0189f
C95 a_15815_855# sigma-delta_0.x1.D 2.42e-20
C96 vpwr a_15706_855# 0.524f
C97 a_15868_1221# a_14791_855# 1.46e-19
C98 a_15141_855# sigma-delta_0.x1.D 0.00353f
C99 a_15596_2320# sigma-delta_0.x1.Q 0.00101f
C100 a_14600_2320# a_14766_3152# 0.00938f
C101 vd sigma-delta_0.x1.D 0.908f
C102 ib buffer_0.a 0.00973f
C103 sensor_0.d sensor_0.c 0.492f
C104 a_15264_2320# a_14932_2320# 0.296f
C105 a_16522_3988# sigma-delta_0.x1.Q 5e-20
C106 ib buffer_0.d 0.766f
C107 out a_15546_5320# 0.00187f
C108 out_buff a_14932_2320# 0.00127f
C109 a_16445_855# sigma-delta_0.in_comp 0.00219f
C110 a_14625_855# sigma-delta_0.in_comp 2.02e-20
C111 a_15380_3988# a_15048_3988# 0.302f
C112 out a_16024_5320# 0.00189f
C113 sigma-delta_0.in_comp sigma-delta_0.in_int 1.13f
C114 out sigma-delta_0.in_int 0.232f
C115 sigma-delta_0.x1.D a_14932_2320# 3.98e-19
C116 a_14625_855# a_15249_1221# 9.73e-19
C117 a_15264_2320# sigma-delta_0.x1.Q 4.28e-19
C118 out_buff buffer_0.b 2.01f
C119 out_sigma a_15706_855# 6.85e-19
C120 a_14791_855# a_15237_855# 2.28e-19
C121 a_15430_3152# sigma-delta_0.x1.Q 2.81e-19
C122 a_15141_855# sigma-delta_0.in_comp 2.02e-20
C123 out_buff buffer_0.a 0.0961f
C124 clk a_15881_829# 2.68e-20
C125 vd out 0.145p
C126 vd sigma-delta_0.in_comp 0.833f
C127 a_15359_1097# sigma-delta_0.x1.Q 0.00111f
C128 a_14766_3152# a_14716_3988# 0.00472f
C129 out_buff buffer_0.d 35.6f
C130 sigma-delta_0.x1.D sigma-delta_0.x1.Q 0.0672f
C131 a_15141_855# a_15249_1221# 0.0572f
C132 a_14625_855# a_15881_829# 0.0436f
C133 a_16445_855# a_15881_829# 0.107f
C134 clk vpwr 0.493f
C135 a_15403_855# vpwr 0.00407f
C136 a_16190_3988# a_16024_5320# 0.00473f
C137 a_16190_3988# sigma-delta_0.in_int 0.358f
C138 out a_16356_5320# 0.00195f
C139 a_15881_829# sigma-delta_0.in_int 0.00137f
C140 a_15046_855# sigma-delta_0.x1.D 0.164f
C141 a_14625_855# vpwr 0.772f
C142 a_16445_855# vpwr 0.2f
C143 sigma-delta_0.in_comp a_14932_2320# 2.76e-19
C144 a_14791_855# a_15596_2320# 1.07e-19
C145 out a_16688_5320# 0.00185f
C146 vd a_16190_3988# 0.00388f
C147 out_buff a_14766_3152# 3.39e-20
C148 vpwr sigma-delta_0.in_int 0.00515f
C149 vd a_15881_829# 0.00172f
C150 a_15264_2320# a_15098_3152# 0.00938f
C151 a_15359_1097# a_15868_1221# 2.6e-19
C152 out buffer_0.b 0.00225f
C153 a_16060_855# sigma-delta_0.x1.D 4.54e-20
C154 a_15815_855# vpwr 7.93e-19
C155 a_16356_5320# a_16190_3988# 0.00536f
C156 a_15868_1221# sigma-delta_0.x1.D 2.11e-20
C157 a_15141_855# vpwr 0.363f
C158 out_buff a_15098_3152# 1.97e-20
C159 a_15430_3152# a_15098_3152# 0.296f
C160 vd vpwr 0.00726f
C161 sigma-delta_0.in_comp sigma-delta_0.x1.Q 0.425f
C162 out_buff a_15214_5320# 5.44e-19
C163 out_sigma clk 0.382f
C164 out buffer_0.a 0.00222f
C165 sigma-delta_0.in_int a_15048_3988# 0.0411f
C166 a_14550_5320# a_14716_3988# 0.00458f
C167 out buffer_0.d 5.5e-19
C168 sigma-delta_0.x1.Q a_15249_1221# 3.66e-19
C169 a_14625_855# out_sigma 0.00261f
C170 out_sigma a_16445_855# 0.0691f
C171 out_buff a_14791_855# 8.29e-20
C172 vd a_15048_3988# 0.00206f
C173 a_15359_1097# a_14791_855# 0.186f
C174 out_buff a_14600_2320# 0.00355f
C175 out_sigma sigma-delta_0.in_int 0.0105f
C176 vts buffer_0.c 0.416f
C177 a_14791_855# sigma-delta_0.x1.D 0.229f
C178 a_15359_1097# a_15237_855# 3.16e-19
C179 sigma-delta_0.x1.Q a_16190_3988# 1.87e-20
C180 a_14766_3152# sigma-delta_0.in_comp 1.21e-19
C181 out_buff a_14550_5320# 0.0535f
C182 a_15881_829# sigma-delta_0.x1.Q 0.142f
C183 a_15237_855# sigma-delta_0.x1.D 8.22e-19
C184 a_15141_855# out_sigma 7.05e-19
C185 vd out_sigma 1.07f
C186 a_15264_2320# a_15596_2320# 0.296f
C187 a_14882_5320# sigma-delta_0.in_int 0.00321f
C188 sigma-delta_0.x1.Q vpwr 0.186f
C189 vd buffer_0.c 0.00573f
C190 sigma-delta_0.in_comp a_15098_3152# 2.91e-19
C191 clk a_15706_855# 6.46e-20
C192 out a_15214_5320# 0.00184f
C193 a_15596_2320# a_15430_3152# 0.00938f
C194 out_buff ib 0.112f
C195 vd a_14882_5320# 0.061f
C196 a_15046_855# vpwr 0.0861f
C197 a_14625_855# a_15706_855# 0.102f
C198 a_16445_855# a_15706_855# 7.05e-19
C199 out_sigma a_14932_2320# 0.0144f
C200 out_buff a_14716_3988# 0.307f
C201 out a_17020_5320# 0.00192f
C202 a_16060_855# a_15881_829# 0.0074f
C203 a_14791_855# sigma-delta_0.in_comp 1.41e-20
C204 a_15380_3988# a_15546_5320# 0.00434f
C205 a_14791_855# a_15249_1221# 0.0346f
C206 out_sigma buffer_0.b 0.0215f
C207 a_15380_3988# sigma-delta_0.in_int 0.339f
C208 a_16060_855# vpwr 0.00312f
C209 out_buff a_15264_2320# 6.31e-19
C210 a_15815_855# a_15706_855# 0.00742f
C211 a_15264_2320# a_15430_3152# 0.00938f
C212 out a_14550_5320# 0.00197f
C213 a_15868_1221# vpwr 9.63e-19
C214 a_15264_2320# a_15359_1097# 1.53e-19
C215 out_sigma sigma-delta_0.x1.Q 0.669f
C216 a_15141_855# a_15706_855# 7.99e-20
C217 vd a_15706_855# 3.52e-19
C218 out_sigma buffer_0.a 0.0182f
C219 buffer_0.b buffer_0.c 0.16f
C220 vd a_15380_3988# 0.00209f
C221 out_buff a_15430_3152# 3.12e-21
C222 out_sigma buffer_0.d 0.00317f
C223 buffer_0.c buffer_0.a 0.199f
C224 a_14791_855# a_15881_829# 0.0426f
C225 out_buff sigma-delta_0.x1.D 1.65e-19
C226 a_15596_2320# sigma-delta_0.in_comp 0.0188f
C227 a_15359_1097# sigma-delta_0.x1.D 6.24e-19
C228 buffer_0.d buffer_0.c 0.0518f
C229 a_15403_855# clk 1.82e-20
C230 a_16522_3988# sigma-delta_0.in_comp 7.16e-19
C231 a_14791_855# vpwr 0.607f
C232 a_15048_3988# a_15098_3152# 0.00472f
C233 a_14625_855# clk 0.274f
C234 a_15214_5320# a_15048_3988# 0.00473f
C235 out_sigma a_14766_3152# 0.00336f
C236 a_15237_855# vpwr 0.00292f
C237 a_14625_855# a_16445_855# 4.71e-20
C238 a_15264_2320# sigma-delta_0.in_comp 4.76e-19
C239 a_16854_3988# sigma-delta_0.in_int 0.0178f
C240 sigma-delta_0.x1.Q a_15706_855# 0.00593f
C241 out_sigma a_15098_3152# 0.00336f
C242 a_16024_5320# a_15546_5320# 0.144f
C243 a_15546_5320# sigma-delta_0.in_int 0.00787f
C244 clk a_15815_855# 1.1e-20
C245 a_16445_855# sigma-delta_0.in_int 0.00209f
C246 a_15141_855# clk 3.26e-19
C247 sigma-delta_0.x1.Q a_15380_3988# 1.43e-21
C248 a_15141_855# a_15403_855# 0.00171f
C249 a_16522_3988# a_16190_3988# 0.312f
C250 out_buff out 0.00558f
C251 a_15430_3152# sigma-delta_0.in_comp 0.297f
C252 a_15359_1097# sigma-delta_0.in_comp 7.49e-21
C253 a_16024_5320# sigma-delta_0.in_int 0.00821f
C254 out a_6126_29386# 0.0171f
C255 a_14625_855# a_15815_855# 2.56e-19
C256 vd a_16854_3988# 0.015f
C257 vd vts 0.94f
C258 vd a_15546_5320# 0.0619f
C259 a_15141_855# a_14625_855# 0.115f
C260 vd a_14625_855# 1.72e-20
C261 out_sigma a_14791_855# 0.00128f
C262 vd a_16445_855# 0.00317f
C263 sigma-delta_0.x1.D sigma-delta_0.in_comp 0.304f
C264 a_15359_1097# a_15249_1221# 0.0977f
C265 out_sigma a_14600_2320# 0.0146f
C266 a_15214_5320# a_14882_5320# 0.303f
C267 vd a_16024_5320# 0.0626f
C268 vd sigma-delta_0.in_int 0.334f
C269 sigma-delta_0.x1.D a_15249_1221# 5.56e-20
C270 out_sigma a_14550_5320# 6.23e-19
C271 out_buff a_16190_3988# 9.87e-22
C272 a_15868_1221# a_15706_855# 0.00645f
C273 a_16356_5320# a_16024_5320# 0.3f
C274 a_16356_5320# sigma-delta_0.in_int 0.00708f
C275 a_14625_855# a_14932_2320# 2.33e-20
C276 a_16688_5320# a_16854_3988# 0.00473f
C277 a_15048_3988# a_14716_3988# 0.296f
C278 a_15264_2320# vpwr 2.29e-19
C279 sigma-delta_0.in_int a_14932_2320# 0.00497f
C280 sigma-delta_0.x1.D a_15881_829# 0.004f
C281 vts buffer_0.b 0.112f
C282 out_buff vpwr 0.00381f
C283 out_sigma a_15596_2320# 0.0144f
C284 a_16688_5320# sigma-delta_0.in_int 0.006f
C285 vts sensor_0.a 0.543f
C286 a_15403_855# sigma-delta_0.x1.Q 9.75e-20
C287 a_14882_5320# a_14550_5320# 0.296f
C288 a_15380_3988# a_15214_5320# 0.00473f
C289 vd a_16356_5320# 0.0637f
C290 a_15359_1097# vpwr 0.378f
C291 clk buffer_0.d 0.0997f
C292 sigma-delta_0.x1.Q a_16854_3988# 0.414f
C293 a_14625_855# sigma-delta_0.x1.Q 9.54e-19
C294 vts buffer_0.a 0.253f
C295 a_16445_855# sigma-delta_0.x1.Q 0.226f
C296 a_14791_855# a_15706_855# 0.125f
C297 sigma-delta_0.x1.D vpwr 0.483f
C298 clk a_15046_855# 3.09e-19
C299 ib buffer_0.c 0.185f
C300 vd a_16688_5320# 0.0633f
C301 vts sensor_0.b 1f
C302 vts buffer_0.d 0.832f
C303 out_buff a_15048_3988# 0.00138f
C304 sigma-delta_0.x1.Q sigma-delta_0.in_int 0.414f
C305 a_14625_855# a_15046_855# 0.0931f
C306 vd buffer_0.b 6.27f
C307 vd sensor_0.a 2.92f
C308 a_15264_2320# out_sigma 0.0144f
C309 a_16060_855# clk 6.32e-21
C310 a_15815_855# sigma-delta_0.x1.Q 1.47e-19
C311 a_16356_5320# a_16688_5320# 0.307f
C312 a_14882_5320# a_14716_3988# 0.00434f
C313 vts sensor_0.c 0.166f
C314 a_15141_855# sigma-delta_0.x1.Q 8.11e-19
C315 vd sigma-delta_0.x1.Q 0.186f
C316 vd buffer_0.a 5.58f
C317 sigma-delta_0.in_comp a_15881_829# 0.00158f
C318 out_buff out_sigma 2.19f
C319 out_sigma a_15430_3152# 0.00336f
C320 out_sigma a_15359_1097# 3.73e-19
C321 vd sensor_0.b 0.0693f
C322 vd buffer_0.d 4.12f
C323 a_15141_855# a_15046_855# 0.0498f
C324 out_sigma sigma-delta_0.x1.D 0.294f
C325 out_buff buffer_0.c 0.0405f
C326 sigma-delta_0.in_comp vpwr 0.00234f
C327 a_14766_3152# sigma-delta_0.in_int 0.399f
C328 vd sensor_0.c 0.804f
C329 clk gnd 2.91f
C330 ib gnd 6.34f
C331 out_buff gnd 14.8f
C332 out gnd 60.4f
C333 out_sigma gnd 18.1f
C334 vpwr gnd 6.13f
C335 vts gnd 19.7f
C336 vd gnd 0.104p
C337 a_16060_855# gnd 0.00223f
C338 a_15815_855# gnd 0.00108f
C339 a_15403_855# gnd 0.00579f
C340 a_15237_855# gnd 0.00863f
C341 a_15868_1221# gnd 3.5e-20
C342 a_15249_1221# gnd 0.00469f
C343 a_15046_855# gnd 0.08f
C344 a_16445_855# gnd 0.213f
C345 a_15706_855# gnd 0.276f
C346 a_15881_829# gnd 0.742f
C347 a_15141_855# gnd 0.282f
C348 a_15359_1097# gnd 0.195f
C349 a_14791_855# gnd 0.334f
C350 sigma-delta_0.x1.D gnd 2.57f
C351 a_14625_855# gnd 0.702f
C352 sigma-delta_0.in_comp gnd 65.9f
C353 a_15596_2320# gnd 0.549f
C354 a_15430_3152# gnd 0.331f
C355 a_15264_2320# gnd 0.349f
C356 a_15098_3152# gnd 0.331f
C357 a_14932_2320# gnd 0.349f
C358 a_14766_3152# gnd 0.331f
C359 a_14600_2320# gnd 0.53f
C360 sigma-delta_0.x1.Q gnd 1.42f
C361 a_17020_5320# gnd 0.52f
C362 a_16854_3988# gnd 0.354f
C363 a_16688_5320# gnd 0.386f
C364 a_16522_3988# gnd 0.361f
C365 a_16356_5320# gnd 0.39f
C366 a_16190_3988# gnd 0.365f
C367 a_16024_5320# gnd 0.444f
C368 sigma-delta_0.in_int gnd 60.9f
C369 a_15546_5320# gnd 0.442f
C370 a_15380_3988# gnd 0.351f
C371 a_15214_5320# gnd 0.38f
C372 a_15048_3988# gnd 0.35f
C373 a_14882_5320# gnd 0.383f
C374 a_14716_3988# gnd 0.35f
C375 a_14550_5320# gnd 0.568f
C376 buffer_0.c gnd 1.15f
C377 buffer_0.b gnd 2.31f
C378 buffer_0.a gnd 2.47f
C379 buffer_0.d gnd 20.2f
C380 sensor_0.b gnd 16.7f
C381 sensor_0.c gnd 0.658f
C382 sensor_0.a gnd 5.59f
C383 sensor_0.d gnd 0.293f
C384 a_6126_29386# gnd 0.593f
C385 out_sigma.t1 gnd 0.0111f
C386 out_sigma.t0 gnd 0.00816f
C387 out_sigma.n0 gnd 0.178f
C388 out_sigma.n1 gnd 0.273f
C389 out_sigma.t2 gnd 0.0241f
C390 out_sigma.n2 gnd 2.11f
C391 out_sigma.n3 gnd 1.36f
C392 out.t0 gnd 0.0079f
C393 out.t3 gnd 13.1f
C394 out.t2 gnd 28.9f
C395 out.t1 gnd 19.8f
C396 out.n0 gnd 10.6f
C397 out.n1 gnd 16.3f
C398 out.n2 gnd 61.4f
C399 vts.t17 gnd 0.1f
C400 vts.t20 gnd 0.00611f
C401 vts.t5 gnd 0.00573f
C402 vts.t3 gnd 0.00573f
C403 vts.n0 gnd 0.0271f
C404 vts.t1 gnd 0.00573f
C405 vts.t16 gnd 0.00573f
C406 vts.n1 gnd 0.0271f
C407 vts.t14 gnd 0.00573f
C408 vts.t12 gnd 0.00573f
C409 vts.n2 gnd 0.0271f
C410 vts.t10 gnd 0.00573f
C411 vts.t8 gnd 0.00573f
C412 vts.n3 gnd 0.0271f
C413 vts.t23 gnd 0.00616f
C414 vts.t21 gnd 0.1f
C415 vts.t24 gnd 0.00603f
C416 vts.n4 gnd 0.12f
C417 vts.n5 gnd 0.0685f
C418 vts.n6 gnd 0.0461f
C419 vts.n7 gnd 0.0538f
C420 vts.n8 gnd 0.0538f
C421 vts.n9 gnd 0.0457f
C422 vts.n10 gnd 0.0683f
C423 vts.n11 gnd 0.0645f
C424 vts.t19 gnd 0.0061f
C425 vts.n12 gnd 0.0548f
C426 vts.n13 gnd 0.00516f
C427 vts.n14 gnd 0.00536f
C428 vts.n15 gnd 0.0344f
C429 vts.n16 gnd 0.0344f
C430 vts.t2 gnd 0.272f
C431 vts.t4 gnd 0.333f
C432 vts.t18 gnd 0.337f
C433 vts.t22 gnd 0.355f
C434 vts.n17 gnd 0.279f
C435 vts.n18 gnd 0.0688f
C436 vts.t0 gnd 0.272f
C437 vts.t15 gnd 0.213f
C438 vts.t7 gnd 0.336f
C439 vts.t9 gnd 0.272f
C440 vts.t11 gnd 0.272f
C441 vts.t13 gnd 0.195f
C442 vts.n19 gnd 0.0653f
C443 vts.n20 gnd 0.0653f
C444 vts.n21 gnd 0.136f
C445 vts.n22 gnd 0.0628f
C446 vts.n23 gnd 0.0628f
C447 vts.n24 gnd 0.0317f
C448 vts.n25 gnd 0.032f
C449 vts.n26 gnd 0.196f
C450 vts.n28 gnd 0.00534f
C451 vts.n29 gnd 0.0103f
C452 vts.n30 gnd 0.00449f
C453 vts.t6 gnd 0.0378f
C454 vts.n31 gnd 0.342f
C455 vts.n32 gnd 8.23e-19
C456 vts.n33 gnd 0.002f
C457 vts.n34 gnd 0.0346f
C458 vts.t25 gnd 0.0138f
C459 vts.n35 gnd 0.669f
C460 vts.n36 gnd 0.833f
C461 buffer_0.d.n0 gnd 0.621f
C462 buffer_0.d.n1 gnd 0.584f
C463 buffer_0.d.t12 gnd 0.274f
C464 buffer_0.d.t13 gnd 0.274f
C465 buffer_0.d.n2 gnd 0.241f
C466 buffer_0.d.t7 gnd 0.274f
C467 buffer_0.d.n3 gnd 0.121f
C468 buffer_0.d.t5 gnd 0.274f
C469 buffer_0.d.n4 gnd 0.149f
C470 buffer_0.d.t9 gnd 33f
C471 buffer_0.d.n5 gnd 0.272f
C472 buffer_0.d.t8 gnd 0.021f
C473 buffer_0.d.t6 gnd 0.021f
C474 buffer_0.d.n6 gnd 0.112f
C475 buffer_0.d.n7 gnd 0.229f
C476 buffer_0.d.t0 gnd 0.701f
C477 buffer_0.d.n8 gnd 0.309f
C478 buffer_0.d.t11 gnd 0.0632f
C479 buffer_0.d.t1 gnd 0.434f
C480 buffer_0.d.t2 gnd 0.701f
C481 buffer_0.d.n9 gnd 0.309f
C482 buffer_0.d.t10 gnd 0.0631f
C483 buffer_0.d.t3 gnd 0.0631f
C484 buffer_0.d.t4 gnd 0.367f
C485 vtd.n0 gnd 0.544f
C486 vtd.n1 gnd 0.544f
C487 vtd.n2 gnd 0.544f
C488 vtd.n3 gnd 0.957f
C489 vtd.n4 gnd 0.174f
C490 vtd.n5 gnd 0.234f
C491 vtd.n6 gnd 0.321f
C492 vtd.t25 gnd 2.06f
C493 vtd.t29 gnd 0.402f
C494 vtd.n7 gnd 1.26f
C495 vtd.t27 gnd 0.401f
C496 vtd.t28 gnd 0.398f
C497 vtd.n8 gnd 0.396f
C498 vtd.t26 gnd 0.398f
C499 vtd.n9 gnd 0.204f
C500 vtd.t24 gnd 0.398f
C501 vtd.t17 gnd 0.0204f
C502 vtd.t21 gnd 0.0115f
C503 vtd.n10 gnd 0.436f
C504 vtd.t18 gnd 0.0115f
C505 vtd.n11 gnd 0.235f
C506 vtd.t22 gnd 0.0114f
C507 vtd.n12 gnd 0.247f
C508 vtd.t19 gnd 0.0114f
C509 vtd.t16 gnd 0.0115f
C510 vtd.t20 gnd 0.0205f
C511 vtd.n13 gnd 0.398f
C512 vtd.t23 gnd 0.0114f
C513 vtd.n14 gnd 0.218f
C514 vtd.n15 gnd 0.322f
C515 vtd.n16 gnd 0.45f
C516 vtd.t5 gnd 0.0239f
C517 vtd.t4 gnd 0.398f
C518 vtd.t12 gnd 0.398f
C519 vtd.t13 gnd 0.0228f
C520 vtd.t7 gnd 0.0228f
C521 vtd.t6 gnd 0.398f
C522 vtd.t0 gnd 0.398f
C523 vtd.t1 gnd 0.0228f
C524 vtd.t9 gnd 0.0228f
C525 vtd.t8 gnd 0.398f
C526 vtd.t14 gnd 0.398f
C527 vtd.t15 gnd 0.0228f
C528 vtd.t11 gnd 0.0228f
C529 vtd.t10 gnd 0.398f
C530 vtd.t2 gnd 0.398f
C531 vtd.t3 gnd 0.0237f
C532 vtd.n17 gnd 0.529f
C533 vtd.n18 gnd 0.339f
C534 vtd.n19 gnd 0.339f
C535 vtd.n20 gnd 0.622f
C536 vd.t74 gnd 21f
C537 vd.t75 gnd 21f
C538 vd.t73 gnd 41.7f
C539 vd.n0 gnd 20.8f
C540 vd.n1 gnd 13.3f
C541 vd.t53 gnd 0.0554f
C542 vd.n2 gnd 17f
C543 vd.n3 gnd 0.0137f
C544 vd.n4 gnd 0.00341f
C545 vd.n5 gnd 0.0104f
C546 vd.n6 gnd 6.52e-19
C547 vd.t17 gnd 0.00767f
C548 vd.n7 gnd 0.00181f
C549 vd.n8 gnd 0.012f
C550 vd.n9 gnd 0.00247f
C551 vd.n10 gnd 0.0138f
C552 vd.n11 gnd 7.05e-19
C553 vd.n12 gnd 0.00505f
C554 vd.n13 gnd 0.0138f
C555 vd.t16 gnd 0.144f
C556 vd.n15 gnd 0.0137f
C557 vd.n16 gnd 0.00505f
C558 vd.n18 gnd 0.139f
C559 vd.n19 gnd 0.0184f
C560 vd.n20 gnd 0.0137f
C561 vd.n21 gnd 0.00562f
C562 vd.n22 gnd 0.00928f
C563 vd.n23 gnd 0.121f
C564 vd.n24 gnd 0.00938f
C565 vd.n25 gnd 0.00574f
C566 vd.n26 gnd 0.0146f
C567 vd.n27 gnd 0.0293f
C568 vd.n28 gnd 0.0148f
C569 vd.n29 gnd 0.0081f
C570 vd.n30 gnd 0.0446f
C571 vd.n31 gnd 0.00316f
C572 vd.n32 gnd 0.00855f
C573 vd.n33 gnd 0.00176f
C574 vd.n34 gnd 0.00229f
C575 vd.n35 gnd 0.00211f
C576 vd.n36 gnd 0.0103f
C577 vd.n37 gnd 0.0136f
C578 vd.n38 gnd 0.218f
C579 vd.n39 gnd 0.0718f
C580 vd.n40 gnd 0.0539f
C581 vd.n41 gnd 0.0798f
C582 vd.n42 gnd 0.585f
C583 vd.t66 gnd -0.0167f
C584 vd.t0 gnd 0.785f
C585 vd.n43 gnd 0.0979f
C586 vd.t37 gnd 0.582f
C587 vd.t52 gnd 0.757f
C588 vd.t35 gnd 0.609f
C589 vd.n44 gnd 0.397f
C590 vd.n45 gnd 0.0646f
C591 vd.n46 gnd 0.0646f
C592 vd.n47 gnd 0.0646f
C593 vd.t28 gnd 0.759f
C594 vd.t29 gnd 0.168f
C595 vd.t31 gnd 0.168f
C596 vd.t33 gnd 0.168f
C597 vd.t42 gnd 0.168f
C598 vd.t39 gnd 0.168f
C599 vd.t41 gnd 0.142f
C600 vd.n48 gnd 0.0678f
C601 vd.n49 gnd 0.0632f
C602 vd.t5 gnd 0.138f
C603 vd.t8 gnd 0.168f
C604 vd.t1 gnd 0.168f
C605 vd.t10 gnd 0.168f
C606 vd.t12 gnd 0.168f
C607 vd.t6 gnd 0.168f
C608 vd.t63 gnd -0.0179f
C609 vd.n50 gnd 0.0798f
C610 vd.t14 gnd 0.595f
C611 vd.n51 gnd 0.398f
C612 vd.t3 gnd 0.598f
C613 vd.t27 gnd 0.755f
C614 vd.n52 gnd 0.623f
C615 vd.n53 gnd 0.0978f
C616 vd.n54 gnd 0.169f
C617 vd.n55 gnd 0.504f
C618 vd.n56 gnd 0.0782f
C619 vd.n57 gnd 0.0782f
C620 vd.n58 gnd 0.0979f
C621 vd.n59 gnd 0.0646f
C622 vd.n60 gnd 0.0792f
C623 vd.n61 gnd 0.0792f
C624 vd.n62 gnd 0.492f
C625 vd.n63 gnd 0.186f
C626 vd.n64 gnd 0.0984f
C627 vd.n65 gnd 0.0715f
C628 vd.n66 gnd 0.0653f
C629 vd.n67 gnd 0.00382f
C630 vd.t40 gnd 0.00255f
C631 vd.t43 gnd 0.00255f
C632 vd.n68 gnd 0.00875f
C633 vd.n69 gnd 0.0086f
C634 vd.t30 gnd 0.00255f
C635 vd.t67 gnd 0.00255f
C636 vd.n70 gnd 0.0116f
C637 vd.t65 gnd 0.0552f
C638 vd.t68 gnd 0.00262f
C639 vd.n71 gnd 0.0813f
C640 vd.n72 gnd 0.022f
C641 vd.t34 gnd 0.00255f
C642 vd.t32 gnd 0.00255f
C643 vd.n73 gnd 0.0143f
C644 vd.n74 gnd 0.0188f
C645 vd.n75 gnd 0.0104f
C646 vd.n76 gnd 0.00127f
C647 vd.n77 gnd 0.0116f
C648 vd.t38 gnd 0.0383f
C649 vd.t36 gnd 0.0383f
C650 vd.n78 gnd 0.324f
C651 vd.n79 gnd 0.271f
C652 vd.t4 gnd 0.0383f
C653 vd.t15 gnd 0.0383f
C654 vd.n80 gnd 0.346f
C655 vd.t62 gnd 0.0552f
C656 vd.n81 gnd 0.0881f
C657 vd.t64 gnd 0.00524f
C658 vd.t7 gnd 0.00255f
C659 vd.n82 gnd 0.0122f
C660 vd.n83 gnd 0.0129f
C661 vd.t13 gnd 0.00255f
C662 vd.t11 gnd 0.00255f
C663 vd.n84 gnd 0.0143f
C664 vd.n85 gnd 0.0196f
C665 vd.t2 gnd 0.00255f
C666 vd.t9 gnd 0.00255f
C667 vd.n86 gnd 0.0105f
C668 vd.n87 gnd 0.0389f
C669 vd.n88 gnd 0.23f
C670 vd.n89 gnd 0.0569f
C671 vd.n90 gnd 0.00405f
C672 vd.n91 gnd 1.23f
C673 vd.t71 gnd 0.00512f
C674 vd.t69 gnd 0.0895f
C675 vd.t72 gnd 0.00512f
C676 vd.t51 gnd 0.00574f
C677 vd.n92 gnd 0.0864f
C678 vd.n93 gnd 0.072f
C679 vd.n94 gnd 0.0921f
C680 vd.n95 gnd 0.0557f
C681 vd.n96 gnd 0.282f
C682 vd.n97 gnd 0.225f
C683 vd.n98 gnd 0.0184f
C684 vd.n99 gnd 0.0184f
C685 vd.t18 gnd 0.091f
C686 vd.t70 gnd 0.0983f
C687 vd.t49 gnd 0.338f
C688 vd.n100 gnd 0.269f
C689 vd.n101 gnd 0.0105f
C690 vd.t48 gnd 0.151f
C691 vd.n102 gnd 0.189f
C692 vd.n103 gnd 0.0138f
C693 vd.n104 gnd 0.0135f
C694 vd.n105 gnd 0.0115f
C695 vd.t58 gnd 0.0896f
C696 vd.t45 gnd 0.00594f
C697 vd.t60 gnd 0.00512f
C698 vd.n106 gnd 0.0838f
C699 vd.n107 gnd 0.0686f
C700 vd.t61 gnd 0.00512f
C701 vd.n108 gnd 0.0727f
C702 vd.n109 gnd 0.00171f
C703 vd.t57 gnd 0.00512f
C704 vd.n110 gnd 0.0297f
C705 vd.t56 gnd 0.00538f
C706 vd.t24 gnd 0.00511f
C707 vd.t26 gnd 0.00511f
C708 vd.n111 gnd 0.0405f
C709 vd.n112 gnd 0.0526f
C710 vd.t54 gnd 0.0894f
C711 vd.n113 gnd 0.0592f
C712 vd.n114 gnd 0.00601f
C713 vd.n115 gnd 0.00276f
C714 vd.n116 gnd 0.0493f
C715 vd.n117 gnd 0.0574f
C716 vd.n118 gnd 0.336f
C717 vd.t55 gnd 0.228f
C718 vd.n119 gnd 0.279f
C719 vd.n120 gnd 0.0217f
C720 vd.n121 gnd 0.0216f
C721 vd.t23 gnd 0.411f
C722 vd.t25 gnd 0.256f
C723 vd.n122 gnd 0.189f
C724 vd.n123 gnd 0.0136f
C725 vd.n124 gnd 0.0147f
C726 vd.n125 gnd 0.115f
C727 vd.n126 gnd 0.139f
C728 vd.t19 gnd 0.0998f
C729 vd.t44 gnd 0.0793f
C730 vd.n127 gnd 0.0818f
C731 vd.n128 gnd 0.0818f
C732 vd.n129 gnd 0.164f
C733 vd.n130 gnd 0.00584f
C734 vd.n131 gnd 0.00582f
C735 vd.t21 gnd 0.244f
C736 vd.n132 gnd 0.28f
C737 vd.n133 gnd 0.0168f
C738 vd.n134 gnd 0.0165f
C739 vd.t20 gnd 0.132f
C740 vd.t22 gnd 0.264f
C741 vd.t59 gnd 0.167f
C742 vd.n135 gnd 0.114f
C743 vd.n136 gnd 0.0111f
C744 vd.n137 gnd 0.0121f
C745 vd.n138 gnd 0.113f
C746 vd.n139 gnd 0.283f
C747 vd.n140 gnd 0.00899f
C748 vd.n141 gnd 0.00888f
C749 vd.t50 gnd 0.189f
C750 vd.t46 gnd 0.186f
C751 vd.t47 gnd 0.286f
C752 vd.n142 gnd 0.189f
C753 vd.n143 gnd 0.0127f
C754 vd.n144 gnd 0.0138f
C755 vd.n145 gnd 0.161f
C756 vd.n146 gnd 0.093f
C757 vd.n147 gnd 0.546f
C758 vd.n148 gnd 5.85f
C759 vd.n149 gnd 4.82f
C760 vd.n150 gnd 0.446f
C761 out_buff.t4 gnd 0.0639f
C762 out_buff.t6 gnd 0.306f
C763 out_buff.t0 gnd 0.0459f
C764 out_buff.n0 gnd 0.169f
C765 out_buff.t5 gnd 0.509f
C766 out_buff.n1 gnd 0.234f
C767 out_buff.n2 gnd 0.0507f
C768 out_buff.t9 gnd 0.263f
C769 out_buff.t1 gnd 0.0459f
C770 out_buff.t8 gnd 0.0459f
C771 out_buff.n3 gnd 0.169f
C772 out_buff.t7 gnd 0.509f
C773 out_buff.n4 gnd 0.233f
C774 out_buff.n5 gnd 0.0508f
C775 out_buff.t11 gnd 0.0103f
C776 out_buff.t10 gnd 38.4f
C777 out_buff.n6 gnd 0.463f
C778 out_buff.t3 gnd 0.0153f
C779 out_buff.t2 gnd 0.0153f
C780 out_buff.n7 gnd 0.11f
C781 out_buff.n8 gnd 0.0705f
C782 out_buff.n9 gnd 0.222f
C783 out_buff.n10 gnd 0.224f
C784 out_buff.n11 gnd 0.493f
C785 out_buff.n12 gnd 1.31f
C786 out_buff.n13 gnd 0.255f
C787 buffer_0.b.n0 gnd 0.0408f
C788 buffer_0.b.n1 gnd 0.0786f
C789 buffer_0.b.t8 gnd 0.0101f
C790 buffer_0.b.t12 gnd 0.0101f
C791 buffer_0.b.n2 gnd 0.0936f
C792 buffer_0.b.t6 gnd 0.0101f
C793 buffer_0.b.t14 gnd 0.0101f
C794 buffer_0.b.n3 gnd 0.0563f
C795 buffer_0.b.n4 gnd 0.0779f
C796 buffer_0.b.n5 gnd 0.0463f
C797 buffer_0.b.t17 gnd 1.68f
C798 buffer_0.b.t16 gnd 1.67f
C799 buffer_0.b.n6 gnd 1.6f
C800 buffer_0.b.t7 gnd 0.126f
C801 buffer_0.b.t11 gnd 0.202f
C802 buffer_0.b.n7 gnd 0.291f
C803 buffer_0.b.t5 gnd 0.202f
C804 buffer_0.b.n8 gnd 0.16f
C805 buffer_0.b.t13 gnd 0.202f
C806 buffer_0.b.n9 gnd 0.16f
C807 buffer_0.b.t9 gnd 0.202f
C808 buffer_0.b.n10 gnd 0.163f
C809 buffer_0.b.t2 gnd 0.202f
C810 buffer_0.b.t4 gnd 0.0104f
C811 buffer_0.b.n11 gnd 0.324f
C812 buffer_0.b.n12 gnd 0.00756f
C813 buffer_0.b.n13 gnd 0.00153f
C814 buffer_0.b.t10 gnd 0.0101f
C815 buffer_0.b.t3 gnd 0.0101f
C816 buffer_0.b.n14 gnd 0.0684f
C817 buffer_0.b.t0 gnd 0.024f
C818 buffer_0.b.t15 gnd 0.0172f
C819 buffer_0.b.t1 gnd 0.0356f
C820 buffer_0.b.n15 gnd 0.224f
C821 buffer_0.b.n16 gnd 0.161f
C822 sensor_0.a.n0 gnd 0.396f
C823 sensor_0.a.n1 gnd 0.413f
C824 sensor_0.a.t15 gnd 0.277f
C825 sensor_0.a.t14 gnd 0.276f
C826 sensor_0.a.n2 gnd 0.293f
C827 sensor_0.a.t12 gnd 0.276f
C828 sensor_0.a.n3 gnd 0.15f
C829 sensor_0.a.t13 gnd 0.276f
C830 sensor_0.a.n4 gnd 0.148f
C831 sensor_0.a.t3 gnd 0.0159f
C832 sensor_0.a.t2 gnd 0.276f
C833 sensor_0.a.t0 gnd 0.276f
C834 sensor_0.a.t1 gnd 0.0177f
C835 sensor_0.a.t11 gnd 0.0141f
C836 sensor_0.a.t8 gnd 0.00791f
C837 sensor_0.a.n5 gnd 0.277f
C838 sensor_0.a.t7 gnd 0.00792f
C839 sensor_0.a.n6 gnd 0.152f
C840 sensor_0.a.t4 gnd 0.00792f
C841 sensor_0.a.n7 gnd 0.19f
C842 sensor_0.a.t6 gnd 0.0141f
C843 sensor_0.a.t10 gnd 0.00791f
C844 sensor_0.a.n8 gnd 0.276f
C845 sensor_0.a.t5 gnd 0.0079f
C846 sensor_0.a.n9 gnd 0.154f
C847 sensor_0.a.t9 gnd 0.00792f
C848 sensor_0.a.n10 gnd 0.19f
C849 sensor_0.a.n11 gnd 0.384f
C850 sensor_0.b.t19 gnd 0.0077f
C851 sensor_0.b.t18 gnd 0.0077f
C852 sensor_0.b.n0 gnd 0.0683f
C853 sensor_0.b.t16 gnd 0.0077f
C854 sensor_0.b.t17 gnd 0.0077f
C855 sensor_0.b.n1 gnd 0.0506f
C856 sensor_0.b.n2 gnd 0.162f
C857 sensor_0.b.t3 gnd 0.00651f
C858 sensor_0.b.t11 gnd 0.00386f
C859 sensor_0.b.n3 gnd 0.139f
C860 sensor_0.b.t5 gnd 0.00385f
C861 sensor_0.b.n4 gnd 0.0928f
C862 sensor_0.b.t13 gnd 0.00385f
C863 sensor_0.b.n5 gnd 0.137f
C864 sensor_0.b.n6 gnd 0.202f
C865 sensor_0.b.t2 gnd 0.134f
C866 sensor_0.b.t10 gnd 0.127f
C867 sensor_0.b.t4 gnd 0.127f
C868 sensor_0.b.t12 gnd 0.0845f
C869 sensor_0.b.t32 gnd 0.134f
C870 sensor_0.b.t24 gnd 0.127f
C871 sensor_0.b.t31 gnd 0.127f
C872 sensor_0.b.t23 gnd 0.0845f
C873 sensor_0.b.t26 gnd 0.134f
C874 sensor_0.b.t34 gnd 0.127f
C875 sensor_0.b.t21 gnd 0.127f
C876 sensor_0.b.t29 gnd 0.0845f
C877 sensor_0.b.t20 gnd 0.134f
C878 sensor_0.b.t27 gnd 0.127f
C879 sensor_0.b.t28 gnd 0.127f
C880 sensor_0.b.t35 gnd 0.0845f
C881 sensor_0.b.t30 gnd 0.134f
C882 sensor_0.b.t22 gnd 0.127f
C883 sensor_0.b.t33 gnd 0.127f
C884 sensor_0.b.t25 gnd 0.0856f
C885 sensor_0.b.n7 gnd 0.119f
C886 sensor_0.b.n8 gnd 0.0626f
C887 sensor_0.b.n9 gnd 0.0626f
C888 sensor_0.b.n10 gnd 0.0626f
C889 sensor_0.b.t0 gnd 0.134f
C890 sensor_0.b.t8 gnd 0.127f
C891 sensor_0.b.t6 gnd 0.127f
C892 sensor_0.b.t14 gnd 0.0845f
C893 sensor_0.b.n11 gnd 0.0519f
C894 sensor_0.b.t1 gnd 0.00705f
C895 sensor_0.b.t9 gnd 0.00386f
C896 sensor_0.b.n12 gnd 0.138f
C897 sensor_0.b.t7 gnd 0.00386f
C898 sensor_0.b.n13 gnd 0.073f
C899 sensor_0.b.t15 gnd 0.00389f
C900 sensor_0.b.n14 gnd 0.0704f
C901 sensor_0.b.n15 gnd 0.0509f
C902 buffer_0.a.n0 gnd 0.146f
C903 buffer_0.a.t11 gnd 0.149f
C904 buffer_0.a.n1 gnd 0.323f
C905 buffer_0.a.t12 gnd 0.014f
C906 buffer_0.a.t4 gnd 0.00689f
C907 buffer_0.a.n2 gnd 0.0272f
C908 buffer_0.a.t3 gnd 0.149f
C909 buffer_0.a.t2 gnd 0.00689f
C910 buffer_0.a.t6 gnd 0.00689f
C911 buffer_0.a.n3 gnd 0.0627f
C912 buffer_0.a.t8 gnd 0.00689f
C913 buffer_0.a.t10 gnd 0.00689f
C914 buffer_0.a.n4 gnd 0.0384f
C915 buffer_0.a.n5 gnd 0.0492f
C916 buffer_0.a.t7 gnd 0.149f
C917 buffer_0.a.t9 gnd 0.149f
C918 buffer_0.a.t1 gnd 0.149f
C919 buffer_0.a.t16 gnd 1.15f
C920 buffer_0.a.t17 gnd 1.15f
C921 buffer_0.a.n6 gnd 0.98f
C922 buffer_0.a.t5 gnd 0.0876f
C923 buffer_0.a.n7 gnd 0.191f
C924 buffer_0.a.n8 gnd 0.0985f
C925 buffer_0.a.n9 gnd 0.0982f
C926 buffer_0.a.n10 gnd 0.026f
C927 buffer_0.a.n11 gnd 0.112f
C928 buffer_0.a.n12 gnd 0.00975f
C929 buffer_0.a.t0 gnd 0.0118f
C930 buffer_0.a.t14 gnd 0.0118f
C931 buffer_0.a.t13 gnd 0.0164f
C932 buffer_0.a.t15 gnd 0.0118f
C933 buffer_0.a.n13 gnd 0.136f
.ends

