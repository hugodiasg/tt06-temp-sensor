VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_hugodg_temp_sensor
  CLASS BLOCK ;
  FOREIGN tt_um_hugodg_temp_sensor ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.000000 ;
    ANTENNADIFFAREA 49.667625 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 30.224998 ;
    ANTENNADIFFAREA 18.850000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.225000 ;
    ANTENNADIFFAREA 12.156000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 120.150 179.800 129.750 196.760 ;
      LAYER nwell ;
        RECT 130.885 179.795 136.215 195.925 ;
        RECT 137.485 175.595 145.815 195.725 ;
        RECT 143.360 168.585 147.060 168.720 ;
        RECT 129.595 161.755 147.060 168.585 ;
      LAYER pwell ;
        RECT 132.260 153.320 143.260 160.220 ;
        RECT 132.260 153.220 137.160 153.320 ;
        RECT 139.360 153.220 143.260 153.320 ;
        RECT 132.260 144.260 143.260 153.220 ;
      LAYER nwell ;
        RECT 143.360 143.620 147.060 161.755 ;
        RECT 129.560 136.820 147.060 143.620 ;
        RECT 125.150 123.960 126.350 125.160 ;
      LAYER pwell ;
        RECT 123.495 123.625 124.175 123.765 ;
        RECT 123.305 123.455 124.175 123.625 ;
        RECT 123.495 119.255 124.175 123.455 ;
      LAYER nwell ;
        RECT 124.695 123.060 126.350 123.960 ;
      LAYER pwell ;
        RECT 123.495 118.325 124.395 119.255 ;
        RECT 123.495 115.605 124.175 118.325 ;
        RECT 123.495 113.250 124.405 115.605 ;
      LAYER nwell ;
        RECT 124.695 113.000 126.300 123.060 ;
      LAYER pwell ;
        RECT 120.670 109.580 123.770 111.690 ;
      LAYER nwell ;
        RECT 124.020 109.580 129.210 111.690 ;
      LAYER pwell ;
        RECT 129.950 109.000 149.050 124.960 ;
      LAYER li1 ;
        RECT 120.330 196.410 129.570 196.580 ;
        RECT 120.330 195.660 120.500 196.410 ;
        RECT 121.420 195.730 122.460 195.900 ;
        RECT 123.510 195.730 124.550 195.900 ;
        RECT 125.600 195.730 126.640 195.900 ;
        RECT 127.690 195.730 128.730 195.900 ;
        RECT 120.330 194.560 120.550 195.660 ;
        RECT 121.080 194.670 121.250 195.670 ;
        RECT 122.630 194.670 122.800 195.670 ;
        RECT 123.170 194.670 123.340 195.670 ;
        RECT 124.720 194.670 124.890 195.670 ;
        RECT 125.260 194.670 125.430 195.670 ;
        RECT 126.810 194.670 126.980 195.670 ;
        RECT 127.350 194.670 127.520 195.670 ;
        RECT 128.900 194.670 129.070 195.670 ;
        RECT 120.330 191.260 120.500 194.560 ;
        RECT 121.420 194.440 122.460 194.610 ;
        RECT 123.510 194.440 124.550 194.610 ;
        RECT 125.600 194.440 126.640 194.610 ;
        RECT 127.690 194.440 128.730 194.610 ;
        RECT 121.420 193.830 122.460 194.000 ;
        RECT 123.510 193.830 124.550 194.000 ;
        RECT 125.600 193.830 126.640 194.000 ;
        RECT 127.690 193.830 128.730 194.000 ;
        RECT 121.080 192.770 121.250 193.770 ;
        RECT 122.630 192.770 122.800 193.770 ;
        RECT 123.170 192.770 123.340 193.770 ;
        RECT 124.720 192.770 124.890 193.770 ;
        RECT 125.260 192.770 125.430 193.770 ;
        RECT 126.810 192.770 126.980 193.770 ;
        RECT 127.350 192.770 127.520 193.770 ;
        RECT 128.900 192.770 129.070 193.770 ;
        RECT 121.420 192.540 122.460 192.710 ;
        RECT 123.510 192.540 124.550 192.710 ;
        RECT 125.600 192.540 126.640 192.710 ;
        RECT 127.690 192.540 128.730 192.710 ;
        RECT 121.420 191.930 122.460 192.100 ;
        RECT 123.510 191.930 124.550 192.100 ;
        RECT 125.600 191.930 126.640 192.100 ;
        RECT 127.690 191.930 128.730 192.100 ;
        RECT 120.330 190.160 120.550 191.260 ;
        RECT 121.080 190.870 121.250 191.870 ;
        RECT 122.630 190.870 122.800 191.870 ;
        RECT 123.170 190.870 123.340 191.870 ;
        RECT 124.720 190.870 124.890 191.870 ;
        RECT 125.260 190.870 125.430 191.870 ;
        RECT 126.810 190.870 126.980 191.870 ;
        RECT 127.350 190.870 127.520 191.870 ;
        RECT 128.900 190.870 129.070 191.870 ;
        RECT 121.420 190.640 122.460 190.810 ;
        RECT 123.510 190.640 124.550 190.810 ;
        RECT 125.600 190.640 126.640 190.810 ;
        RECT 127.690 190.640 128.730 190.810 ;
        RECT 120.330 186.660 120.500 190.160 ;
        RECT 121.420 190.030 122.460 190.200 ;
        RECT 123.510 190.030 124.550 190.200 ;
        RECT 125.600 190.030 126.640 190.200 ;
        RECT 127.690 190.030 128.730 190.200 ;
        RECT 121.080 188.970 121.250 189.970 ;
        RECT 122.630 188.970 122.800 189.970 ;
        RECT 123.170 188.970 123.340 189.970 ;
        RECT 124.720 188.970 124.890 189.970 ;
        RECT 125.260 188.970 125.430 189.970 ;
        RECT 126.810 188.970 126.980 189.970 ;
        RECT 127.350 188.970 127.520 189.970 ;
        RECT 128.900 188.970 129.070 189.970 ;
        RECT 121.420 188.740 122.460 188.910 ;
        RECT 123.510 188.740 124.550 188.910 ;
        RECT 125.600 188.740 126.640 188.910 ;
        RECT 127.690 188.740 128.730 188.910 ;
        RECT 121.420 188.130 122.460 188.300 ;
        RECT 123.510 188.130 124.550 188.300 ;
        RECT 125.600 188.130 126.640 188.300 ;
        RECT 127.690 188.130 128.730 188.300 ;
        RECT 121.080 187.070 121.250 188.070 ;
        RECT 122.630 187.070 122.800 188.070 ;
        RECT 123.170 187.070 123.340 188.070 ;
        RECT 124.720 187.070 124.890 188.070 ;
        RECT 125.260 187.070 125.430 188.070 ;
        RECT 126.810 187.070 126.980 188.070 ;
        RECT 127.350 187.070 127.520 188.070 ;
        RECT 128.900 187.070 129.070 188.070 ;
        RECT 121.420 186.840 122.460 187.010 ;
        RECT 123.510 186.840 124.550 187.010 ;
        RECT 125.600 186.840 126.640 187.010 ;
        RECT 127.690 186.840 128.730 187.010 ;
        RECT 120.330 185.560 120.550 186.660 ;
        RECT 121.420 186.230 122.460 186.400 ;
        RECT 123.510 186.230 124.550 186.400 ;
        RECT 125.600 186.230 126.640 186.400 ;
        RECT 127.690 186.230 128.730 186.400 ;
        RECT 120.330 182.460 120.500 185.560 ;
        RECT 121.080 185.170 121.250 186.170 ;
        RECT 122.630 185.170 122.800 186.170 ;
        RECT 123.170 185.170 123.340 186.170 ;
        RECT 124.720 185.170 124.890 186.170 ;
        RECT 125.260 185.170 125.430 186.170 ;
        RECT 126.810 185.170 126.980 186.170 ;
        RECT 127.350 185.170 127.520 186.170 ;
        RECT 128.900 185.170 129.070 186.170 ;
        RECT 121.420 184.940 122.460 185.110 ;
        RECT 123.510 184.940 124.550 185.110 ;
        RECT 125.600 184.940 126.640 185.110 ;
        RECT 127.690 184.940 128.730 185.110 ;
        RECT 121.420 184.330 122.460 184.500 ;
        RECT 123.510 184.330 124.550 184.500 ;
        RECT 125.600 184.330 126.640 184.500 ;
        RECT 127.690 184.330 128.730 184.500 ;
        RECT 121.080 183.270 121.250 184.270 ;
        RECT 122.630 183.270 122.800 184.270 ;
        RECT 123.170 183.270 123.340 184.270 ;
        RECT 124.720 183.270 124.890 184.270 ;
        RECT 125.260 183.270 125.430 184.270 ;
        RECT 126.810 183.270 126.980 184.270 ;
        RECT 127.350 183.270 127.520 184.270 ;
        RECT 128.900 183.270 129.070 184.270 ;
        RECT 121.420 183.040 122.460 183.210 ;
        RECT 123.510 183.040 124.550 183.210 ;
        RECT 125.600 183.040 126.640 183.210 ;
        RECT 127.690 183.040 128.730 183.210 ;
        RECT 120.330 181.360 120.550 182.460 ;
        RECT 121.420 182.430 122.460 182.600 ;
        RECT 123.510 182.430 124.550 182.600 ;
        RECT 125.600 182.430 126.640 182.600 ;
        RECT 127.690 182.430 128.730 182.600 ;
        RECT 121.080 181.370 121.250 182.370 ;
        RECT 122.630 181.370 122.800 182.370 ;
        RECT 123.170 181.370 123.340 182.370 ;
        RECT 124.720 181.370 124.890 182.370 ;
        RECT 125.260 181.370 125.430 182.370 ;
        RECT 126.810 181.370 126.980 182.370 ;
        RECT 127.350 181.370 127.520 182.370 ;
        RECT 128.900 181.370 129.070 182.370 ;
        RECT 120.330 180.150 120.500 181.360 ;
        RECT 121.420 181.140 122.460 181.310 ;
        RECT 123.510 181.140 124.550 181.310 ;
        RECT 125.600 181.140 126.640 181.310 ;
        RECT 127.690 181.140 128.730 181.310 ;
        RECT 129.400 180.150 129.570 196.410 ;
        RECT 120.330 179.980 129.570 180.150 ;
        RECT 131.065 195.575 136.035 195.745 ;
        RECT 131.065 180.145 131.235 195.575 ;
        RECT 132.630 194.750 134.670 194.920 ;
        RECT 132.245 193.690 132.415 194.690 ;
        RECT 134.885 193.690 135.055 194.690 ;
        RECT 132.630 193.460 134.670 193.630 ;
        RECT 132.630 192.850 134.670 193.020 ;
        RECT 132.245 191.790 132.415 192.790 ;
        RECT 134.885 191.790 135.055 192.790 ;
        RECT 132.630 191.560 134.670 191.730 ;
        RECT 132.245 190.500 132.415 191.500 ;
        RECT 134.885 190.500 135.055 191.500 ;
        RECT 132.630 190.270 134.670 190.440 ;
        RECT 132.245 189.210 132.415 190.210 ;
        RECT 134.885 189.210 135.055 190.210 ;
        RECT 132.630 188.980 134.670 189.150 ;
        RECT 132.245 187.920 132.415 188.920 ;
        RECT 134.885 187.920 135.055 188.920 ;
        RECT 132.630 187.690 134.670 187.860 ;
        RECT 132.245 186.630 132.415 187.630 ;
        RECT 134.885 186.630 135.055 187.630 ;
        RECT 132.630 186.400 134.670 186.570 ;
        RECT 132.245 185.340 132.415 186.340 ;
        RECT 134.885 185.340 135.055 186.340 ;
        RECT 132.630 185.110 134.670 185.280 ;
        RECT 132.245 184.050 132.415 185.050 ;
        RECT 134.885 184.050 135.055 185.050 ;
        RECT 132.630 183.820 134.670 183.990 ;
        RECT 132.245 182.760 132.415 183.760 ;
        RECT 134.885 182.760 135.055 183.760 ;
        RECT 132.630 182.530 134.670 182.700 ;
        RECT 132.630 181.950 134.670 182.120 ;
        RECT 132.245 180.890 132.415 181.890 ;
        RECT 134.885 180.890 135.055 181.890 ;
        RECT 132.630 180.660 134.670 180.830 ;
        RECT 134.050 180.145 134.550 180.360 ;
        RECT 135.865 180.145 136.035 195.575 ;
        RECT 131.065 179.975 136.035 180.145 ;
        RECT 137.665 195.375 145.635 195.545 ;
        RECT 134.050 179.960 134.550 179.975 ;
        RECT 137.665 175.945 137.835 195.375 ;
        RECT 138.830 194.650 140.870 194.820 ;
        RECT 138.445 193.590 138.615 194.590 ;
        RECT 141.085 193.590 141.255 194.590 ;
        RECT 138.830 193.360 140.870 193.530 ;
        RECT 138.830 192.750 140.870 192.920 ;
        RECT 138.445 191.690 138.615 192.690 ;
        RECT 141.085 191.690 141.255 192.690 ;
        RECT 145.465 192.560 145.635 195.375 ;
        RECT 145.450 191.760 145.650 192.560 ;
        RECT 138.830 191.460 140.870 191.630 ;
        RECT 138.445 190.400 138.615 191.400 ;
        RECT 141.085 190.400 141.255 191.400 ;
        RECT 138.830 190.170 140.870 190.340 ;
        RECT 138.830 189.550 140.870 189.720 ;
        RECT 138.445 188.490 138.615 189.490 ;
        RECT 141.085 188.490 141.255 189.490 ;
        RECT 138.830 188.260 140.870 188.430 ;
        RECT 138.445 187.200 138.615 188.200 ;
        RECT 141.085 187.200 141.255 188.200 ;
        RECT 142.230 187.750 144.270 187.920 ;
        RECT 138.830 186.970 140.870 187.140 ;
        RECT 138.445 185.910 138.615 186.910 ;
        RECT 141.085 185.910 141.255 186.910 ;
        RECT 141.845 186.690 142.015 187.690 ;
        RECT 144.485 186.690 144.655 187.690 ;
        RECT 145.465 186.960 145.635 191.760 ;
        RECT 142.230 186.460 144.270 186.630 ;
        RECT 145.450 186.160 145.650 186.960 ;
        RECT 142.230 185.850 144.270 186.020 ;
        RECT 138.830 185.680 140.870 185.850 ;
        RECT 138.445 184.620 138.615 185.620 ;
        RECT 141.085 184.620 141.255 185.620 ;
        RECT 141.845 184.790 142.015 185.790 ;
        RECT 144.485 184.790 144.655 185.790 ;
        RECT 142.230 184.560 144.270 184.730 ;
        RECT 138.830 184.390 140.870 184.560 ;
        RECT 142.230 183.950 144.270 184.120 ;
        RECT 138.830 183.750 140.870 183.920 ;
        RECT 138.445 182.690 138.615 183.690 ;
        RECT 141.085 182.690 141.255 183.690 ;
        RECT 138.830 182.460 140.870 182.630 ;
        RECT 138.445 181.400 138.615 182.400 ;
        RECT 141.085 181.400 141.255 182.400 ;
        RECT 138.830 181.170 140.870 181.340 ;
        RECT 138.445 180.110 138.615 181.110 ;
        RECT 141.085 180.110 141.255 181.110 ;
        RECT 138.830 179.880 140.870 180.050 ;
        RECT 138.445 178.820 138.615 179.820 ;
        RECT 141.085 178.820 141.255 179.820 ;
        RECT 141.845 178.890 142.015 183.890 ;
        RECT 144.485 178.890 144.655 183.890 ;
        RECT 145.465 183.060 145.635 186.160 ;
        RECT 145.450 182.260 145.650 183.060 ;
        RECT 138.830 178.590 140.870 178.760 ;
        RECT 142.230 178.660 144.270 178.830 ;
        RECT 145.465 178.460 145.635 182.260 ;
        RECT 138.830 177.950 140.870 178.120 ;
        RECT 142.230 178.050 144.270 178.220 ;
        RECT 138.445 176.890 138.615 177.890 ;
        RECT 141.085 176.890 141.255 177.890 ;
        RECT 141.845 176.990 142.015 177.990 ;
        RECT 144.485 176.990 144.655 177.990 ;
        RECT 145.450 177.660 145.650 178.460 ;
        RECT 138.830 176.660 140.870 176.830 ;
        RECT 142.230 176.760 144.270 176.930 ;
        RECT 145.465 175.945 145.635 177.660 ;
        RECT 137.665 175.775 145.635 175.945 ;
        RECT 129.775 168.235 146.845 168.405 ;
        RECT 129.775 162.105 129.945 168.235 ;
        RECT 143.575 168.220 143.745 168.235 ;
        RECT 130.740 167.710 145.780 167.880 ;
        RECT 130.355 166.650 130.525 167.650 ;
        RECT 145.995 166.650 146.165 167.650 ;
        RECT 130.740 166.420 145.780 166.590 ;
        RECT 130.355 165.360 130.525 166.360 ;
        RECT 145.995 165.360 146.165 166.360 ;
        RECT 130.740 165.130 145.780 165.300 ;
        RECT 130.355 164.070 130.525 165.070 ;
        RECT 145.995 164.070 146.165 165.070 ;
        RECT 130.740 163.840 145.780 164.010 ;
        RECT 130.355 162.780 130.525 163.780 ;
        RECT 145.995 162.780 146.165 163.780 ;
        RECT 130.740 162.550 145.780 162.720 ;
        RECT 143.175 162.105 143.745 162.120 ;
        RECT 129.775 162.020 143.745 162.105 ;
        RECT 129.775 161.935 143.760 162.020 ;
        RECT 143.560 160.720 143.760 161.935 ;
        RECT 144.740 161.910 145.780 162.080 ;
        RECT 144.355 160.850 144.525 161.850 ;
        RECT 145.995 160.850 146.165 161.850 ;
        RECT 146.675 161.405 146.845 168.235 ;
        RECT 146.660 161.235 146.845 161.405 ;
        RECT 132.440 159.870 143.180 160.040 ;
        RECT 132.440 156.220 132.610 159.870 ;
        RECT 137.780 158.490 138.820 158.660 ;
        RECT 137.440 157.430 137.610 158.430 ;
        RECT 138.990 157.430 139.160 158.430 ;
        RECT 137.780 157.200 138.820 157.370 ;
        RECT 132.360 155.720 132.760 156.220 ;
        RECT 137.440 156.140 137.610 157.140 ;
        RECT 138.990 156.140 139.160 157.140 ;
        RECT 137.780 155.910 138.820 156.080 ;
        RECT 132.440 149.120 132.610 155.720 ;
        RECT 137.440 154.850 137.610 155.850 ;
        RECT 138.990 154.850 139.160 155.850 ;
        RECT 137.780 154.620 138.820 154.790 ;
        RECT 137.440 153.560 137.610 154.560 ;
        RECT 138.990 153.560 139.160 154.560 ;
        RECT 137.780 153.330 138.820 153.500 ;
        RECT 140.540 153.070 140.710 153.400 ;
        RECT 140.880 153.390 142.420 153.560 ;
        RECT 140.880 152.910 142.420 153.080 ;
        RECT 133.480 152.690 138.520 152.860 ;
        RECT 133.140 151.630 133.310 152.630 ;
        RECT 138.690 151.630 138.860 152.630 ;
        RECT 140.540 152.110 140.710 152.440 ;
        RECT 140.880 152.430 142.420 152.600 ;
        RECT 142.590 152.590 142.760 152.920 ;
        RECT 140.880 151.950 142.420 152.120 ;
        RECT 133.480 151.400 138.520 151.570 ;
        RECT 140.880 151.470 142.420 151.640 ;
        RECT 142.590 151.630 142.760 151.960 ;
        RECT 133.140 150.340 133.310 151.340 ;
        RECT 138.690 150.340 138.860 151.340 ;
        RECT 133.480 150.110 138.520 150.280 ;
        RECT 132.360 148.620 132.760 149.120 ;
        RECT 133.140 149.050 133.310 150.050 ;
        RECT 138.690 149.050 138.860 150.050 ;
        RECT 133.480 148.820 138.520 148.990 ;
        RECT 132.440 144.610 132.610 148.620 ;
        RECT 133.140 147.760 133.310 148.760 ;
        RECT 138.690 147.760 138.860 148.760 ;
        RECT 133.480 147.530 138.520 147.700 ;
        RECT 133.140 146.470 133.310 147.470 ;
        RECT 138.690 146.470 138.860 147.470 ;
        RECT 133.480 146.240 138.520 146.410 ;
        RECT 133.140 145.180 133.310 146.180 ;
        RECT 138.690 145.180 138.860 146.180 ;
        RECT 133.480 144.950 138.520 145.120 ;
        RECT 143.010 144.610 143.180 159.870 ;
        RECT 132.440 144.440 143.180 144.610 ;
        RECT 143.575 143.405 143.745 160.720 ;
        RECT 144.740 160.620 145.780 160.790 ;
        RECT 144.355 159.560 144.525 160.560 ;
        RECT 145.995 159.560 146.165 160.560 ;
        RECT 144.740 159.330 145.780 159.500 ;
        RECT 144.355 158.270 144.525 159.270 ;
        RECT 145.995 158.270 146.165 159.270 ;
        RECT 144.740 158.040 145.780 158.210 ;
        RECT 144.355 156.980 144.525 157.980 ;
        RECT 145.995 156.980 146.165 157.980 ;
        RECT 144.740 156.750 145.780 156.920 ;
        RECT 144.355 155.690 144.525 156.690 ;
        RECT 145.995 155.690 146.165 156.690 ;
        RECT 144.740 155.460 145.780 155.630 ;
        RECT 144.355 154.400 144.525 155.400 ;
        RECT 145.995 154.400 146.165 155.400 ;
        RECT 146.675 155.320 146.845 161.235 ;
        RECT 144.740 154.170 145.780 154.340 ;
        RECT 144.355 153.110 144.525 154.110 ;
        RECT 145.995 153.110 146.165 154.110 ;
        RECT 144.740 152.880 145.780 153.050 ;
        RECT 144.740 152.310 145.780 152.480 ;
        RECT 144.355 151.230 144.525 152.250 ;
        RECT 145.995 151.250 146.165 152.250 ;
        RECT 144.740 151.020 145.780 151.190 ;
        RECT 144.355 149.940 144.525 150.960 ;
        RECT 145.995 149.960 146.165 150.960 ;
        RECT 146.660 150.120 146.860 155.320 ;
        RECT 144.740 149.730 145.780 149.900 ;
        RECT 144.355 148.650 144.525 149.670 ;
        RECT 145.995 148.670 146.165 149.670 ;
        RECT 144.740 148.440 145.780 148.610 ;
        RECT 144.355 147.360 144.525 148.380 ;
        RECT 145.995 147.380 146.165 148.380 ;
        RECT 144.740 147.150 145.780 147.320 ;
        RECT 144.355 146.070 144.525 147.090 ;
        RECT 145.995 146.090 146.165 147.090 ;
        RECT 144.740 145.860 145.780 146.030 ;
        RECT 144.355 144.800 144.525 145.800 ;
        RECT 145.995 144.800 146.165 145.800 ;
        RECT 144.740 144.570 145.780 144.740 ;
        RECT 144.355 143.490 144.525 144.510 ;
        RECT 145.995 143.510 146.165 144.510 ;
        RECT 146.675 143.905 146.845 150.120 ;
        RECT 146.660 143.735 146.845 143.905 ;
        RECT 129.775 143.235 143.760 143.405 ;
        RECT 144.740 143.280 145.780 143.450 ;
        RECT 129.775 137.205 129.945 143.235 ;
        RECT 130.740 142.710 145.780 142.880 ;
        RECT 130.355 141.650 130.525 142.650 ;
        RECT 145.995 141.650 146.165 142.650 ;
        RECT 130.740 141.420 145.780 141.590 ;
        RECT 130.355 140.360 130.525 141.360 ;
        RECT 145.995 140.360 146.165 141.360 ;
        RECT 130.740 140.130 145.780 140.300 ;
        RECT 130.355 139.070 130.525 140.070 ;
        RECT 145.995 139.070 146.165 140.070 ;
        RECT 130.740 138.840 145.780 139.010 ;
        RECT 130.355 137.780 130.525 138.780 ;
        RECT 145.995 137.780 146.165 138.780 ;
        RECT 130.740 137.550 145.780 137.720 ;
        RECT 146.675 137.520 146.845 143.735 ;
        RECT 143.575 137.205 143.745 137.220 ;
        RECT 146.660 137.205 146.860 137.520 ;
        RECT 129.775 137.035 146.860 137.205 ;
        RECT 146.660 137.020 146.860 137.035 ;
        RECT 125.450 124.160 125.900 124.660 ;
        RECT 130.130 124.610 148.870 124.780 ;
        RECT 123.305 123.255 123.475 123.770 ;
        RECT 123.735 123.425 124.195 123.680 ;
        RECT 123.305 122.925 123.855 123.255 ;
        RECT 124.025 123.160 124.195 123.425 ;
        RECT 124.365 123.330 125.015 123.680 ;
        RECT 125.185 123.425 125.855 123.680 ;
        RECT 125.185 123.160 125.355 123.425 ;
        RECT 126.025 123.255 126.195 123.770 ;
        RECT 124.025 122.930 125.355 123.160 ;
        RECT 125.525 122.925 126.195 123.255 ;
        RECT 123.305 122.225 123.475 122.925 ;
        RECT 123.735 122.585 125.855 122.755 ;
        RECT 125.055 122.355 125.840 122.415 ;
        RECT 123.305 121.895 123.835 122.225 ;
        RECT 124.005 122.090 125.840 122.355 ;
        RECT 124.005 121.895 125.055 122.090 ;
        RECT 126.025 121.920 126.195 122.925 ;
        RECT 123.305 119.295 123.475 121.895 ;
        RECT 123.695 121.555 125.395 121.725 ;
        RECT 125.565 121.670 126.195 121.920 ;
        RECT 123.695 121.230 123.865 121.555 ;
        RECT 125.225 121.500 125.395 121.555 ;
        RECT 124.155 121.035 124.775 121.385 ;
        RECT 125.225 121.330 125.855 121.500 ;
        RECT 125.525 121.250 125.855 121.330 ;
        RECT 123.695 120.340 123.865 121.025 ;
        RECT 124.965 120.865 125.355 121.160 ;
        RECT 124.155 120.695 125.355 120.865 ;
        RECT 124.155 120.510 124.375 120.695 ;
        RECT 125.525 120.525 125.855 121.035 ;
        RECT 124.575 120.355 125.855 120.525 ;
        RECT 124.575 120.340 124.745 120.355 ;
        RECT 123.695 120.170 124.745 120.340 ;
        RECT 123.305 118.965 123.935 119.295 ;
        RECT 124.155 119.175 124.405 119.965 ;
        RECT 124.575 119.005 124.745 120.170 ;
        RECT 125.255 120.015 125.765 120.185 ;
        RECT 123.305 117.065 123.475 118.965 ;
        RECT 124.395 118.835 124.745 119.005 ;
        RECT 123.665 118.665 124.225 118.755 ;
        RECT 124.915 118.665 125.085 119.995 ;
        RECT 125.255 119.280 125.425 120.015 ;
        RECT 126.025 119.780 126.195 121.670 ;
        RECT 125.595 119.450 126.195 119.780 ;
        RECT 125.255 119.110 125.765 119.280 ;
        RECT 126.025 118.815 126.195 119.450 ;
        RECT 123.665 118.495 125.395 118.665 ;
        RECT 123.665 118.405 123.835 118.495 ;
        RECT 123.645 117.405 123.925 118.185 ;
        RECT 124.095 118.095 125.055 118.305 ;
        RECT 125.225 118.275 125.395 118.495 ;
        RECT 125.565 118.445 126.195 118.815 ;
        RECT 125.225 118.105 125.855 118.275 ;
        RECT 124.095 117.575 124.715 117.925 ;
        RECT 124.885 117.800 125.055 118.095 ;
        RECT 124.885 117.630 125.345 117.800 ;
        RECT 123.645 117.235 124.875 117.405 ;
        RECT 125.045 117.340 125.345 117.630 ;
        RECT 124.705 117.170 124.875 117.235 ;
        RECT 125.515 117.170 125.855 117.870 ;
        RECT 123.305 116.875 123.915 117.065 ;
        RECT 123.305 115.435 123.475 116.875 ;
        RECT 124.085 116.845 124.535 117.065 ;
        RECT 124.705 117.000 125.855 117.170 ;
        RECT 124.085 116.705 124.255 116.845 ;
        RECT 123.685 116.535 124.255 116.705 ;
        RECT 123.685 115.955 123.855 116.535 ;
        RECT 124.425 116.365 124.795 116.665 ;
        RECT 124.025 116.125 124.795 116.365 ;
        RECT 123.685 115.780 124.685 115.955 ;
        RECT 124.965 115.950 125.135 117.000 ;
        RECT 126.025 116.830 126.195 118.445 ;
        RECT 125.565 116.580 126.195 116.830 ;
        RECT 125.305 116.240 125.765 116.410 ;
        RECT 125.305 115.780 125.475 116.240 ;
        RECT 126.025 116.060 126.195 116.580 ;
        RECT 123.685 115.635 125.475 115.780 ;
        RECT 124.210 115.630 125.475 115.635 ;
        RECT 124.385 115.610 125.475 115.630 ;
        RECT 123.305 115.265 124.160 115.435 ;
        RECT 124.385 115.335 124.715 115.610 ;
        RECT 125.645 115.340 126.195 116.060 ;
        RECT 123.305 114.010 123.475 115.265 ;
        RECT 124.845 115.095 125.855 115.170 ;
        RECT 123.665 114.765 125.855 115.095 ;
        RECT 123.850 114.760 124.150 114.765 ;
        RECT 123.735 114.325 125.815 114.575 ;
        RECT 124.385 114.245 125.815 114.325 ;
        RECT 123.305 113.840 124.070 114.010 ;
        RECT 123.305 113.190 123.475 113.840 ;
        RECT 124.385 113.715 124.715 114.245 ;
        RECT 126.025 114.010 126.195 115.340 ;
        RECT 124.885 113.840 126.195 114.010 ;
        RECT 123.655 113.545 124.185 113.590 ;
        RECT 124.835 113.545 125.715 113.590 ;
        RECT 123.655 113.335 125.715 113.545 ;
        RECT 124.450 113.310 124.650 113.335 ;
        RECT 126.025 113.190 126.195 113.840 ;
        RECT 130.130 116.660 130.300 124.610 ;
        RECT 130.950 123.410 133.110 123.760 ;
        RECT 135.110 123.410 137.270 123.760 ;
        RECT 139.290 123.660 141.450 124.010 ;
        RECT 145.950 123.660 148.110 124.010 ;
        RECT 130.950 122.580 133.110 122.930 ;
        RECT 135.110 122.580 137.270 122.930 ;
        RECT 139.290 122.830 141.450 123.180 ;
        RECT 145.950 122.830 148.110 123.180 ;
        RECT 130.950 121.750 133.110 122.100 ;
        RECT 135.110 121.750 137.270 122.100 ;
        RECT 139.290 122.000 141.450 122.350 ;
        RECT 145.950 122.000 148.110 122.350 ;
        RECT 130.950 120.920 133.110 121.270 ;
        RECT 135.110 120.920 137.270 121.270 ;
        RECT 139.290 121.170 141.450 121.520 ;
        RECT 145.950 121.170 148.110 121.520 ;
        RECT 130.950 120.090 133.110 120.440 ;
        RECT 135.110 120.090 137.270 120.440 ;
        RECT 139.290 120.340 141.450 120.690 ;
        RECT 145.950 120.340 148.110 120.690 ;
        RECT 130.950 119.260 133.110 119.610 ;
        RECT 135.110 119.260 137.270 119.610 ;
        RECT 139.290 119.510 141.450 119.860 ;
        RECT 145.950 119.510 148.110 119.860 ;
        RECT 130.950 118.430 133.110 118.780 ;
        RECT 135.110 118.430 137.270 118.780 ;
        RECT 139.290 118.680 141.450 119.030 ;
        RECT 145.950 118.680 148.110 119.030 ;
        RECT 130.950 117.600 133.110 117.950 ;
        RECT 135.110 117.600 137.270 117.950 ;
        RECT 139.290 117.850 141.450 118.200 ;
        RECT 145.950 117.850 148.110 118.200 ;
        RECT 130.130 116.060 130.350 116.660 ;
        RECT 139.290 116.290 141.450 116.640 ;
        RECT 145.950 116.290 148.110 116.640 ;
        RECT 120.850 111.340 123.590 111.510 ;
        RECT 120.850 109.930 121.020 111.340 ;
        RECT 121.360 110.470 121.530 110.800 ;
        RECT 121.700 110.770 122.740 110.940 ;
        RECT 121.700 110.330 122.740 110.500 ;
        RECT 122.910 110.470 123.080 110.800 ;
        RECT 121.750 109.930 122.550 109.960 ;
        RECT 123.420 109.930 123.590 111.340 ;
        RECT 120.850 109.760 123.590 109.930 ;
        RECT 124.200 111.340 129.030 111.510 ;
        RECT 124.200 109.930 124.370 111.340 ;
        RECT 124.710 110.470 124.880 110.800 ;
        RECT 125.095 110.770 128.135 110.940 ;
        RECT 125.095 110.330 128.135 110.500 ;
        RECT 128.350 110.470 128.520 110.800 ;
        RECT 125.250 109.930 128.050 109.960 ;
        RECT 128.860 109.930 129.030 111.340 ;
        RECT 124.200 109.760 129.030 109.930 ;
        RECT 130.130 109.350 130.300 116.060 ;
        RECT 139.290 115.460 141.450 115.810 ;
        RECT 145.950 115.460 148.110 115.810 ;
        RECT 139.290 114.630 141.450 114.980 ;
        RECT 145.950 114.630 148.110 114.980 ;
        RECT 139.290 113.800 141.450 114.150 ;
        RECT 145.950 113.800 148.110 114.150 ;
        RECT 139.290 112.970 141.450 113.320 ;
        RECT 145.950 112.970 148.110 113.320 ;
        RECT 139.290 112.140 141.450 112.490 ;
        RECT 145.950 112.140 148.110 112.490 ;
        RECT 139.290 111.310 141.450 111.660 ;
        RECT 145.950 111.310 148.110 111.660 ;
        RECT 139.290 110.480 141.450 110.830 ;
        RECT 145.950 110.480 148.110 110.830 ;
        RECT 148.700 109.350 148.870 124.610 ;
        RECT 130.130 109.180 148.870 109.350 ;
      LAYER mcon ;
        RECT 121.500 195.730 122.380 195.900 ;
        RECT 123.590 195.730 124.470 195.900 ;
        RECT 125.680 195.730 126.560 195.900 ;
        RECT 127.770 195.730 128.650 195.900 ;
        RECT 120.350 194.560 120.550 195.660 ;
        RECT 121.080 194.750 121.250 195.590 ;
        RECT 122.630 194.750 122.800 195.590 ;
        RECT 123.170 194.750 123.340 195.590 ;
        RECT 124.720 194.750 124.890 195.590 ;
        RECT 125.260 194.750 125.430 195.590 ;
        RECT 126.810 194.750 126.980 195.590 ;
        RECT 127.350 194.750 127.520 195.590 ;
        RECT 128.900 194.750 129.070 195.590 ;
        RECT 121.500 194.440 122.380 194.610 ;
        RECT 123.590 194.440 124.470 194.610 ;
        RECT 125.680 194.440 126.560 194.610 ;
        RECT 127.770 194.440 128.650 194.610 ;
        RECT 121.500 193.830 122.380 194.000 ;
        RECT 123.590 193.830 124.470 194.000 ;
        RECT 125.680 193.830 126.560 194.000 ;
        RECT 127.770 193.830 128.650 194.000 ;
        RECT 121.080 192.850 121.250 193.690 ;
        RECT 122.630 192.850 122.800 193.690 ;
        RECT 123.170 192.850 123.340 193.690 ;
        RECT 124.720 192.850 124.890 193.690 ;
        RECT 125.260 192.850 125.430 193.690 ;
        RECT 126.810 192.850 126.980 193.690 ;
        RECT 127.350 192.850 127.520 193.690 ;
        RECT 128.900 192.850 129.070 193.690 ;
        RECT 121.500 192.540 122.380 192.710 ;
        RECT 123.590 192.540 124.470 192.710 ;
        RECT 125.680 192.540 126.560 192.710 ;
        RECT 127.770 192.540 128.650 192.710 ;
        RECT 121.500 191.930 122.380 192.100 ;
        RECT 123.590 191.930 124.470 192.100 ;
        RECT 125.680 191.930 126.560 192.100 ;
        RECT 127.770 191.930 128.650 192.100 ;
        RECT 120.350 190.160 120.550 191.260 ;
        RECT 121.080 190.950 121.250 191.790 ;
        RECT 122.630 190.950 122.800 191.790 ;
        RECT 123.170 190.950 123.340 191.790 ;
        RECT 124.720 190.950 124.890 191.790 ;
        RECT 125.260 190.950 125.430 191.790 ;
        RECT 126.810 190.950 126.980 191.790 ;
        RECT 127.350 190.950 127.520 191.790 ;
        RECT 128.900 190.950 129.070 191.790 ;
        RECT 121.500 190.640 122.380 190.810 ;
        RECT 123.590 190.640 124.470 190.810 ;
        RECT 125.680 190.640 126.560 190.810 ;
        RECT 127.770 190.640 128.650 190.810 ;
        RECT 121.500 190.030 122.380 190.200 ;
        RECT 123.590 190.030 124.470 190.200 ;
        RECT 125.680 190.030 126.560 190.200 ;
        RECT 127.770 190.030 128.650 190.200 ;
        RECT 121.080 189.050 121.250 189.890 ;
        RECT 122.630 189.050 122.800 189.890 ;
        RECT 123.170 189.050 123.340 189.890 ;
        RECT 124.720 189.050 124.890 189.890 ;
        RECT 125.260 189.050 125.430 189.890 ;
        RECT 126.810 189.050 126.980 189.890 ;
        RECT 127.350 189.050 127.520 189.890 ;
        RECT 128.900 189.050 129.070 189.890 ;
        RECT 121.500 188.740 122.380 188.910 ;
        RECT 123.590 188.740 124.470 188.910 ;
        RECT 125.680 188.740 126.560 188.910 ;
        RECT 127.770 188.740 128.650 188.910 ;
        RECT 121.500 188.130 122.380 188.300 ;
        RECT 123.590 188.130 124.470 188.300 ;
        RECT 125.680 188.130 126.560 188.300 ;
        RECT 127.770 188.130 128.650 188.300 ;
        RECT 121.080 187.150 121.250 187.990 ;
        RECT 122.630 187.150 122.800 187.990 ;
        RECT 123.170 187.150 123.340 187.990 ;
        RECT 124.720 187.150 124.890 187.990 ;
        RECT 125.260 187.150 125.430 187.990 ;
        RECT 126.810 187.150 126.980 187.990 ;
        RECT 127.350 187.150 127.520 187.990 ;
        RECT 128.900 187.150 129.070 187.990 ;
        RECT 121.500 186.840 122.380 187.010 ;
        RECT 123.590 186.840 124.470 187.010 ;
        RECT 125.680 186.840 126.560 187.010 ;
        RECT 127.770 186.840 128.650 187.010 ;
        RECT 120.350 185.560 120.550 186.660 ;
        RECT 121.500 186.230 122.380 186.400 ;
        RECT 123.590 186.230 124.470 186.400 ;
        RECT 125.680 186.230 126.560 186.400 ;
        RECT 127.770 186.230 128.650 186.400 ;
        RECT 121.080 185.250 121.250 186.090 ;
        RECT 122.630 185.250 122.800 186.090 ;
        RECT 123.170 185.250 123.340 186.090 ;
        RECT 124.720 185.250 124.890 186.090 ;
        RECT 125.260 185.250 125.430 186.090 ;
        RECT 126.810 185.250 126.980 186.090 ;
        RECT 127.350 185.250 127.520 186.090 ;
        RECT 128.900 185.250 129.070 186.090 ;
        RECT 121.500 184.940 122.380 185.110 ;
        RECT 123.590 184.940 124.470 185.110 ;
        RECT 125.680 184.940 126.560 185.110 ;
        RECT 127.770 184.940 128.650 185.110 ;
        RECT 121.500 184.330 122.380 184.500 ;
        RECT 123.590 184.330 124.470 184.500 ;
        RECT 125.680 184.330 126.560 184.500 ;
        RECT 127.770 184.330 128.650 184.500 ;
        RECT 121.080 183.350 121.250 184.190 ;
        RECT 122.630 183.350 122.800 184.190 ;
        RECT 123.170 183.350 123.340 184.190 ;
        RECT 124.720 183.350 124.890 184.190 ;
        RECT 125.260 183.350 125.430 184.190 ;
        RECT 126.810 183.350 126.980 184.190 ;
        RECT 127.350 183.350 127.520 184.190 ;
        RECT 128.900 183.350 129.070 184.190 ;
        RECT 121.500 183.040 122.380 183.210 ;
        RECT 123.590 183.040 124.470 183.210 ;
        RECT 125.680 183.040 126.560 183.210 ;
        RECT 127.770 183.040 128.650 183.210 ;
        RECT 120.350 181.360 120.550 182.460 ;
        RECT 121.500 182.430 122.380 182.600 ;
        RECT 123.590 182.430 124.470 182.600 ;
        RECT 125.680 182.430 126.560 182.600 ;
        RECT 127.770 182.430 128.650 182.600 ;
        RECT 121.080 181.450 121.250 182.290 ;
        RECT 122.630 181.450 122.800 182.290 ;
        RECT 123.170 181.450 123.340 182.290 ;
        RECT 124.720 181.450 124.890 182.290 ;
        RECT 125.260 181.450 125.430 182.290 ;
        RECT 126.810 181.450 126.980 182.290 ;
        RECT 127.350 181.450 127.520 182.290 ;
        RECT 128.900 181.450 129.070 182.290 ;
        RECT 121.500 181.140 122.380 181.310 ;
        RECT 123.590 181.140 124.470 181.310 ;
        RECT 125.680 181.140 126.560 181.310 ;
        RECT 127.770 181.140 128.650 181.310 ;
        RECT 133.565 194.750 134.505 194.920 ;
        RECT 132.245 193.770 132.415 194.610 ;
        RECT 134.885 193.770 135.055 194.610 ;
        RECT 133.565 193.460 134.505 193.630 ;
        RECT 132.795 192.850 133.735 193.020 ;
        RECT 132.245 191.870 132.415 192.710 ;
        RECT 134.885 191.870 135.055 192.710 ;
        RECT 133.565 191.560 134.505 191.730 ;
        RECT 132.245 190.580 132.415 191.420 ;
        RECT 134.885 190.580 135.055 191.420 ;
        RECT 132.795 190.270 133.735 190.440 ;
        RECT 132.245 189.290 132.415 190.130 ;
        RECT 134.885 189.290 135.055 190.130 ;
        RECT 133.565 188.980 134.505 189.150 ;
        RECT 132.245 188.000 132.415 188.840 ;
        RECT 134.885 188.000 135.055 188.840 ;
        RECT 132.795 187.690 133.735 187.860 ;
        RECT 132.245 186.710 132.415 187.550 ;
        RECT 134.885 186.710 135.055 187.550 ;
        RECT 133.565 186.400 134.505 186.570 ;
        RECT 132.245 185.420 132.415 186.260 ;
        RECT 134.885 185.420 135.055 186.260 ;
        RECT 132.795 185.110 133.735 185.280 ;
        RECT 132.245 184.130 132.415 184.970 ;
        RECT 134.885 184.130 135.055 184.970 ;
        RECT 133.565 183.820 134.505 183.990 ;
        RECT 132.245 182.840 132.415 183.680 ;
        RECT 134.885 182.840 135.055 183.680 ;
        RECT 132.795 182.530 133.735 182.700 ;
        RECT 133.565 181.950 134.505 182.120 ;
        RECT 132.245 180.970 132.415 181.810 ;
        RECT 134.885 180.970 135.055 181.810 ;
        RECT 133.565 180.660 134.505 180.830 ;
        RECT 139.765 194.650 140.705 194.820 ;
        RECT 138.445 193.670 138.615 194.510 ;
        RECT 141.085 193.670 141.255 194.510 ;
        RECT 139.765 193.360 140.705 193.530 ;
        RECT 138.995 192.750 139.935 192.920 ;
        RECT 138.445 191.770 138.615 192.610 ;
        RECT 141.085 191.770 141.255 192.610 ;
        RECT 145.450 191.760 145.650 192.560 ;
        RECT 139.765 191.460 140.705 191.630 ;
        RECT 138.445 190.480 138.615 191.320 ;
        RECT 141.085 190.480 141.255 191.320 ;
        RECT 138.995 190.170 139.935 190.340 ;
        RECT 138.995 189.550 139.935 189.720 ;
        RECT 138.445 188.570 138.615 189.410 ;
        RECT 141.085 188.570 141.255 189.410 ;
        RECT 139.765 188.260 140.705 188.430 ;
        RECT 138.445 187.280 138.615 188.120 ;
        RECT 141.085 187.280 141.255 188.120 ;
        RECT 143.165 187.750 144.105 187.920 ;
        RECT 138.995 186.970 139.935 187.140 ;
        RECT 138.445 185.990 138.615 186.830 ;
        RECT 141.085 185.990 141.255 186.830 ;
        RECT 141.845 186.770 142.015 187.610 ;
        RECT 144.485 186.770 144.655 187.610 ;
        RECT 143.165 186.460 144.105 186.630 ;
        RECT 145.450 186.160 145.650 186.960 ;
        RECT 142.310 185.850 144.190 186.020 ;
        RECT 139.765 185.680 140.705 185.850 ;
        RECT 138.445 184.700 138.615 185.540 ;
        RECT 141.085 184.700 141.255 185.540 ;
        RECT 141.845 184.870 142.015 185.710 ;
        RECT 144.485 184.870 144.655 185.710 ;
        RECT 142.310 184.560 144.190 184.730 ;
        RECT 138.995 184.390 139.935 184.560 ;
        RECT 142.310 183.950 144.190 184.120 ;
        RECT 138.995 183.750 139.935 183.920 ;
        RECT 138.445 182.770 138.615 183.610 ;
        RECT 141.085 182.770 141.255 183.610 ;
        RECT 139.765 182.460 140.705 182.630 ;
        RECT 138.445 181.480 138.615 182.320 ;
        RECT 141.085 181.480 141.255 182.320 ;
        RECT 138.995 181.170 139.935 181.340 ;
        RECT 138.445 180.190 138.615 181.030 ;
        RECT 141.085 180.190 141.255 181.030 ;
        RECT 139.765 179.880 140.705 180.050 ;
        RECT 138.445 178.900 138.615 179.740 ;
        RECT 141.085 178.900 141.255 179.740 ;
        RECT 141.845 178.970 142.015 183.810 ;
        RECT 144.485 178.970 144.655 183.810 ;
        RECT 145.450 182.260 145.650 183.060 ;
        RECT 138.995 178.590 139.935 178.760 ;
        RECT 142.310 178.660 144.190 178.830 ;
        RECT 138.995 177.950 139.935 178.120 ;
        RECT 143.165 178.050 144.105 178.220 ;
        RECT 138.445 176.970 138.615 177.810 ;
        RECT 141.085 176.970 141.255 177.810 ;
        RECT 141.845 177.070 142.015 177.910 ;
        RECT 144.485 177.070 144.655 177.910 ;
        RECT 145.450 177.660 145.650 178.460 ;
        RECT 138.995 176.660 139.935 176.830 ;
        RECT 143.165 176.760 144.105 176.930 ;
        RECT 138.175 167.710 145.615 167.880 ;
        RECT 130.355 166.730 130.525 167.570 ;
        RECT 130.905 166.420 138.345 166.590 ;
        RECT 145.995 165.440 146.165 166.280 ;
        RECT 138.175 165.130 145.615 165.300 ;
        RECT 145.995 164.150 146.165 164.990 ;
        RECT 130.905 163.840 138.345 164.010 ;
        RECT 130.355 162.860 130.525 163.700 ;
        RECT 138.175 162.550 145.615 162.720 ;
        RECT 144.905 161.910 145.345 162.080 ;
        RECT 144.355 160.930 144.525 161.770 ;
        RECT 137.945 158.490 138.385 158.660 ;
        RECT 137.440 157.510 137.610 158.350 ;
        RECT 138.990 157.510 139.160 158.350 ;
        RECT 138.215 157.200 138.655 157.370 ;
        RECT 137.440 156.220 137.610 157.060 ;
        RECT 132.360 155.720 132.760 156.220 ;
        RECT 138.990 156.220 139.160 157.060 ;
        RECT 137.945 155.910 138.385 156.080 ;
        RECT 137.440 154.930 137.610 155.770 ;
        RECT 138.990 154.930 139.160 155.770 ;
        RECT 138.215 154.620 138.655 154.790 ;
        RECT 137.440 153.640 137.610 154.480 ;
        RECT 138.990 153.640 139.160 154.480 ;
        RECT 137.945 153.330 138.385 153.500 ;
        RECT 141.045 153.390 141.735 153.560 ;
        RECT 140.540 153.150 140.710 153.320 ;
        RECT 141.565 152.910 142.255 153.080 ;
        RECT 135.915 152.690 138.355 152.860 ;
        RECT 142.590 152.670 142.760 152.840 ;
        RECT 133.140 151.710 133.310 152.550 ;
        RECT 138.690 151.710 138.860 152.550 ;
        RECT 141.045 152.430 141.735 152.600 ;
        RECT 140.540 152.190 140.710 152.360 ;
        RECT 141.565 151.950 142.255 152.120 ;
        RECT 142.590 151.710 142.760 151.880 ;
        RECT 133.645 151.400 136.085 151.570 ;
        RECT 141.045 151.470 141.735 151.640 ;
        RECT 133.140 150.420 133.310 151.260 ;
        RECT 138.690 150.420 138.860 151.260 ;
        RECT 135.915 150.110 138.355 150.280 ;
        RECT 133.140 149.130 133.310 149.970 ;
        RECT 132.360 148.620 132.760 149.120 ;
        RECT 138.690 149.130 138.860 149.970 ;
        RECT 133.645 148.820 136.085 148.990 ;
        RECT 133.140 147.840 133.310 148.680 ;
        RECT 138.690 147.840 138.860 148.680 ;
        RECT 135.915 147.530 138.355 147.700 ;
        RECT 133.140 146.550 133.310 147.390 ;
        RECT 138.690 146.550 138.860 147.390 ;
        RECT 133.645 146.240 136.085 146.410 ;
        RECT 133.140 145.260 133.310 146.100 ;
        RECT 138.690 145.260 138.860 146.100 ;
        RECT 135.915 144.950 138.355 145.120 ;
        RECT 145.175 160.620 145.615 160.790 ;
        RECT 144.355 159.640 144.525 160.480 ;
        RECT 145.995 159.640 146.165 160.480 ;
        RECT 144.905 159.330 145.345 159.500 ;
        RECT 144.355 158.350 144.525 159.190 ;
        RECT 145.175 158.040 145.615 158.210 ;
        RECT 144.355 157.060 144.525 157.900 ;
        RECT 144.905 156.750 145.345 156.920 ;
        RECT 144.355 155.770 144.525 156.610 ;
        RECT 145.175 155.460 145.615 155.630 ;
        RECT 144.355 154.480 144.525 155.320 ;
        RECT 144.905 154.170 145.345 154.340 ;
        RECT 144.355 153.190 144.525 154.030 ;
        RECT 145.175 152.880 145.615 153.050 ;
        RECT 144.905 152.310 145.345 152.480 ;
        RECT 145.175 151.020 145.615 151.190 ;
        RECT 146.660 150.120 146.860 155.320 ;
        RECT 144.905 149.730 145.345 149.900 ;
        RECT 145.175 148.440 145.615 148.610 ;
        RECT 144.905 147.150 145.345 147.320 ;
        RECT 145.175 145.860 145.615 146.030 ;
        RECT 144.355 144.880 144.525 145.720 ;
        RECT 145.995 144.880 146.165 145.720 ;
        RECT 144.905 144.570 145.345 144.740 ;
        RECT 145.175 143.280 145.615 143.450 ;
        RECT 138.175 142.710 145.615 142.880 ;
        RECT 130.355 141.730 130.525 142.570 ;
        RECT 130.905 141.420 138.345 141.590 ;
        RECT 145.995 140.440 146.165 141.280 ;
        RECT 138.175 140.130 145.615 140.300 ;
        RECT 145.995 139.150 146.165 139.990 ;
        RECT 130.905 138.840 138.345 139.010 ;
        RECT 130.355 137.860 130.525 138.700 ;
        RECT 138.175 137.550 145.615 137.720 ;
        RECT 125.600 124.260 125.850 124.610 ;
        RECT 123.305 123.455 123.475 123.625 ;
        RECT 123.305 122.995 123.475 123.165 ;
        RECT 124.450 123.460 124.750 123.660 ;
        RECT 126.025 123.455 126.195 123.625 ;
        RECT 124.495 122.990 124.665 123.160 ;
        RECT 126.025 122.995 126.195 123.165 ;
        RECT 123.305 122.535 123.475 122.705 ;
        RECT 125.175 122.585 125.345 122.755 ;
        RECT 126.025 122.535 126.195 122.705 ;
        RECT 123.305 122.075 123.475 122.245 ;
        RECT 124.100 121.960 124.300 122.260 ;
        RECT 126.025 122.075 126.195 122.245 ;
        RECT 123.305 121.615 123.475 121.785 ;
        RECT 123.305 121.155 123.475 121.325 ;
        RECT 126.025 121.615 126.195 121.785 ;
        RECT 124.495 121.155 124.665 121.325 ;
        RECT 123.305 120.695 123.475 120.865 ;
        RECT 123.305 120.235 123.475 120.405 ;
        RECT 126.025 121.155 126.195 121.325 ;
        RECT 125.175 120.695 125.345 120.865 ;
        RECT 126.025 120.695 126.195 120.865 ;
        RECT 126.025 120.235 126.195 120.405 ;
        RECT 123.305 119.775 123.475 119.945 ;
        RECT 123.305 119.315 123.475 119.485 ;
        RECT 124.155 119.795 124.325 119.965 ;
        RECT 124.155 119.435 124.325 119.605 ;
        RECT 123.305 118.855 123.475 119.025 ;
        RECT 123.305 118.395 123.475 118.565 ;
        RECT 126.025 119.775 126.195 119.945 ;
        RECT 126.025 119.315 126.195 119.485 ;
        RECT 126.025 118.855 126.195 119.025 ;
        RECT 123.305 117.935 123.475 118.105 ;
        RECT 123.305 117.475 123.475 117.645 ;
        RECT 126.025 118.395 126.195 118.565 ;
        RECT 124.495 117.575 124.665 117.745 ;
        RECT 126.025 117.935 126.195 118.105 ;
        RECT 125.175 117.575 125.345 117.745 ;
        RECT 123.305 117.015 123.475 117.185 ;
        RECT 123.305 116.555 123.475 116.725 ;
        RECT 126.025 117.475 126.195 117.645 ;
        RECT 126.025 117.015 126.195 117.185 ;
        RECT 123.305 116.095 123.475 116.265 ;
        RECT 123.305 115.635 123.475 115.805 ;
        RECT 124.470 116.495 124.640 116.665 ;
        RECT 124.155 116.195 124.325 116.365 ;
        RECT 126.025 116.555 126.195 116.725 ;
        RECT 126.025 116.095 126.195 116.265 ;
        RECT 126.025 115.635 126.195 115.805 ;
        RECT 123.305 115.175 123.475 115.345 ;
        RECT 126.025 115.175 126.195 115.345 ;
        RECT 123.305 114.715 123.475 114.885 ;
        RECT 126.025 114.715 126.195 114.885 ;
        RECT 123.305 114.255 123.475 114.425 ;
        RECT 126.025 114.255 126.195 114.425 ;
        RECT 123.305 113.795 123.475 113.965 ;
        RECT 126.025 113.795 126.195 113.965 ;
        RECT 123.305 113.335 123.475 113.505 ;
        RECT 126.025 113.335 126.195 113.505 ;
        RECT 131.040 123.490 133.025 123.680 ;
        RECT 135.195 123.490 137.180 123.680 ;
        RECT 139.380 123.740 141.365 123.930 ;
        RECT 146.035 123.740 148.020 123.930 ;
        RECT 131.040 122.660 133.025 122.850 ;
        RECT 135.195 122.660 137.180 122.850 ;
        RECT 139.380 122.910 141.365 123.100 ;
        RECT 146.035 122.910 148.020 123.100 ;
        RECT 131.040 121.830 133.025 122.020 ;
        RECT 135.195 121.830 137.180 122.020 ;
        RECT 139.380 122.080 141.365 122.270 ;
        RECT 146.035 122.080 148.020 122.270 ;
        RECT 131.040 121.000 133.025 121.190 ;
        RECT 135.195 121.000 137.180 121.190 ;
        RECT 139.380 121.250 141.365 121.440 ;
        RECT 146.035 121.250 148.020 121.440 ;
        RECT 131.040 120.170 133.025 120.360 ;
        RECT 135.195 120.170 137.180 120.360 ;
        RECT 139.380 120.420 141.365 120.610 ;
        RECT 146.035 120.420 148.020 120.610 ;
        RECT 131.040 119.340 133.025 119.530 ;
        RECT 135.195 119.340 137.180 119.530 ;
        RECT 139.380 119.590 141.365 119.780 ;
        RECT 146.035 119.590 148.020 119.780 ;
        RECT 131.040 118.510 133.025 118.700 ;
        RECT 135.195 118.510 137.180 118.700 ;
        RECT 139.380 118.760 141.365 118.950 ;
        RECT 146.035 118.760 148.020 118.950 ;
        RECT 131.040 117.680 133.025 117.870 ;
        RECT 135.195 117.680 137.180 117.870 ;
        RECT 139.380 117.930 141.365 118.120 ;
        RECT 146.035 117.930 148.020 118.120 ;
        RECT 139.380 116.370 141.365 116.560 ;
        RECT 146.035 116.370 148.020 116.560 ;
        RECT 121.780 110.770 122.660 110.940 ;
        RECT 121.360 110.550 121.530 110.720 ;
        RECT 122.910 110.550 123.080 110.720 ;
        RECT 121.780 110.330 122.660 110.500 ;
        RECT 121.750 109.760 122.550 109.960 ;
        RECT 125.175 110.770 128.055 110.940 ;
        RECT 124.710 110.550 124.880 110.720 ;
        RECT 128.350 110.550 128.520 110.720 ;
        RECT 125.175 110.330 128.055 110.500 ;
        RECT 125.250 109.760 128.050 109.960 ;
        RECT 139.380 115.540 141.365 115.730 ;
        RECT 146.035 115.540 148.020 115.730 ;
        RECT 139.380 114.710 141.365 114.900 ;
        RECT 146.035 114.710 148.020 114.900 ;
        RECT 139.380 113.880 141.365 114.070 ;
        RECT 146.035 113.880 148.020 114.070 ;
        RECT 139.380 113.050 141.365 113.240 ;
        RECT 146.035 113.050 148.020 113.240 ;
        RECT 139.380 112.220 141.365 112.410 ;
        RECT 146.035 112.220 148.020 112.410 ;
        RECT 139.380 111.390 141.365 111.580 ;
        RECT 146.035 111.390 148.020 111.580 ;
        RECT 139.380 110.560 141.365 110.750 ;
        RECT 146.035 110.560 148.020 110.750 ;
      LAYER met1 ;
        RECT 109.570 196.470 110.570 197.070 ;
        RECT 107.870 174.970 108.370 175.020 ;
        RECT 107.870 174.960 108.470 174.970 ;
        RECT 106.450 173.970 108.470 174.960 ;
        RECT 106.450 173.960 108.370 173.970 ;
        RECT 107.870 173.920 108.370 173.960 ;
        RECT 107.850 171.970 108.550 172.010 ;
        RECT 106.470 170.970 108.570 171.970 ;
        RECT 107.850 170.910 108.550 170.970 ;
        RECT 106.470 130.370 108.570 131.370 ;
        RECT 106.470 128.270 107.470 128.470 ;
        RECT 106.470 127.470 108.470 128.270 ;
        RECT 107.870 126.670 108.470 126.720 ;
        RECT 106.470 125.870 108.470 126.670 ;
        RECT 106.470 125.670 107.470 125.870 ;
        RECT 107.870 125.820 108.470 125.870 ;
        RECT 106.470 125.270 107.470 125.370 ;
        RECT 106.470 124.370 108.570 125.270 ;
        RECT 107.470 124.270 108.570 124.370 ;
        RECT 109.170 116.270 111.370 196.470 ;
        RECT 119.350 194.360 129.200 195.960 ;
        RECT 134.050 194.950 134.550 194.960 ;
        RECT 133.505 194.860 134.565 194.950 ;
        RECT 133.505 194.720 135.150 194.860 ;
        RECT 140.450 194.850 140.850 195.210 ;
        RECT 119.350 191.320 120.400 194.360 ;
        RECT 121.500 194.030 122.400 194.110 ;
        RECT 123.600 194.030 124.500 194.110 ;
        RECT 125.600 194.030 126.600 194.110 ;
        RECT 127.800 194.030 128.700 194.110 ;
        RECT 121.440 193.800 122.440 194.030 ;
        RECT 123.530 193.800 124.530 194.030 ;
        RECT 125.600 193.800 126.620 194.030 ;
        RECT 127.710 193.800 128.710 194.030 ;
        RECT 121.050 192.790 121.280 193.750 ;
        RECT 121.500 193.710 122.400 193.800 ;
        RECT 122.600 193.460 122.830 193.750 ;
        RECT 123.140 193.460 123.370 193.750 ;
        RECT 123.600 193.710 124.500 193.800 ;
        RECT 122.600 192.960 123.370 193.460 ;
        RECT 122.600 192.790 122.830 192.960 ;
        RECT 123.140 192.790 123.370 192.960 ;
        RECT 124.690 193.460 124.920 193.750 ;
        RECT 125.230 193.460 125.460 193.750 ;
        RECT 125.600 193.710 126.600 193.800 ;
        RECT 124.690 192.960 125.460 193.460 ;
        RECT 124.690 192.790 124.920 192.960 ;
        RECT 125.230 192.790 125.460 192.960 ;
        RECT 126.780 193.460 127.010 193.750 ;
        RECT 127.320 193.460 127.550 193.750 ;
        RECT 127.800 193.710 128.700 193.800 ;
        RECT 128.950 193.750 129.150 193.760 ;
        RECT 126.780 192.960 127.550 193.460 ;
        RECT 126.780 192.790 127.010 192.960 ;
        RECT 127.320 192.790 127.550 192.960 ;
        RECT 128.870 192.790 129.150 193.750 ;
        RECT 121.440 192.510 122.440 192.740 ;
        RECT 123.530 192.710 124.530 192.740 ;
        RECT 125.620 192.710 126.620 192.740 ;
        RECT 127.710 192.710 128.710 192.740 ;
        RECT 123.500 192.510 124.530 192.710 ;
        RECT 125.600 192.510 126.620 192.710 ;
        RECT 127.700 192.510 128.710 192.710 ;
        RECT 121.500 192.130 122.400 192.510 ;
        RECT 123.500 192.130 124.500 192.510 ;
        RECT 125.600 192.130 126.600 192.510 ;
        RECT 127.700 192.130 128.700 192.510 ;
        RECT 121.440 191.900 122.440 192.130 ;
        RECT 123.500 191.910 124.530 192.130 ;
        RECT 125.600 191.910 126.620 192.130 ;
        RECT 127.700 191.910 128.710 192.130 ;
        RECT 123.530 191.900 124.530 191.910 ;
        RECT 125.620 191.900 126.620 191.910 ;
        RECT 127.710 191.900 128.710 191.910 ;
        RECT 128.950 191.850 129.150 192.790 ;
        RECT 119.350 190.100 120.580 191.320 ;
        RECT 121.050 190.890 121.280 191.850 ;
        RECT 122.600 191.660 122.830 191.850 ;
        RECT 123.140 191.660 123.370 191.850 ;
        RECT 122.600 191.160 123.370 191.660 ;
        RECT 121.500 190.840 122.400 190.910 ;
        RECT 122.600 190.890 122.830 191.160 ;
        RECT 123.140 190.890 123.370 191.160 ;
        RECT 124.690 191.660 124.920 191.850 ;
        RECT 125.230 191.660 125.460 191.850 ;
        RECT 126.780 191.660 127.010 191.850 ;
        RECT 127.320 191.660 127.550 191.850 ;
        RECT 124.690 191.160 125.460 191.660 ;
        RECT 126.750 191.160 127.550 191.660 ;
        RECT 123.600 190.840 124.500 190.910 ;
        RECT 124.690 190.890 124.920 191.160 ;
        RECT 125.230 190.890 125.460 191.160 ;
        RECT 125.700 190.840 126.600 190.910 ;
        RECT 126.780 190.890 127.010 191.160 ;
        RECT 127.320 190.890 127.550 191.160 ;
        RECT 127.800 190.840 128.700 190.910 ;
        RECT 128.870 190.890 129.150 191.850 ;
        RECT 121.440 190.610 122.440 190.840 ;
        RECT 123.530 190.610 124.530 190.840 ;
        RECT 125.620 190.610 126.620 190.840 ;
        RECT 127.710 190.610 128.710 190.840 ;
        RECT 121.500 190.510 122.400 190.610 ;
        RECT 123.600 190.510 124.500 190.610 ;
        RECT 125.700 190.510 126.600 190.610 ;
        RECT 127.800 190.510 128.700 190.610 ;
        RECT 121.500 190.230 122.300 190.310 ;
        RECT 123.600 190.230 124.400 190.310 ;
        RECT 125.700 190.230 126.500 190.310 ;
        RECT 127.800 190.230 128.600 190.310 ;
        RECT 119.350 186.720 120.400 190.100 ;
        RECT 121.440 190.000 122.440 190.230 ;
        RECT 123.530 190.000 124.530 190.230 ;
        RECT 125.620 190.000 126.620 190.230 ;
        RECT 127.710 190.000 128.710 190.230 ;
        RECT 121.050 188.990 121.280 189.950 ;
        RECT 121.500 189.910 122.300 190.000 ;
        RECT 122.600 189.760 122.830 189.950 ;
        RECT 123.140 189.760 123.370 189.950 ;
        RECT 123.600 189.910 124.400 190.000 ;
        RECT 122.600 189.260 123.370 189.760 ;
        RECT 122.600 188.990 122.830 189.260 ;
        RECT 123.140 188.990 123.370 189.260 ;
        RECT 124.690 189.760 124.920 189.950 ;
        RECT 125.230 189.760 125.460 189.950 ;
        RECT 125.700 189.910 126.500 190.000 ;
        RECT 126.780 189.760 127.010 189.950 ;
        RECT 127.320 189.760 127.550 189.950 ;
        RECT 127.800 189.910 128.600 190.000 ;
        RECT 128.950 189.950 129.150 190.890 ;
        RECT 130.550 190.510 130.950 194.110 ;
        RECT 132.215 193.710 132.445 194.670 ;
        RECT 134.050 193.660 135.150 194.720 ;
        RECT 139.705 194.620 140.850 194.850 ;
        RECT 133.505 193.560 135.150 193.660 ;
        RECT 138.415 193.610 138.645 194.570 ;
        RECT 140.450 194.560 140.850 194.620 ;
        RECT 145.850 195.160 146.350 195.210 ;
        RECT 141.055 194.560 141.285 194.570 ;
        RECT 140.450 193.610 141.285 194.560 ;
        RECT 140.450 193.560 141.250 193.610 ;
        RECT 133.505 193.430 134.565 193.560 ;
        RECT 132.150 193.050 133.350 193.060 ;
        RECT 132.150 192.820 133.795 193.050 ;
        RECT 132.150 190.470 133.350 192.820 ;
        RECT 134.050 191.760 134.550 193.430 ;
        RECT 139.705 193.330 140.850 193.560 ;
        RECT 138.550 192.950 139.450 192.960 ;
        RECT 134.855 191.810 135.085 192.770 ;
        RECT 138.550 192.720 139.995 192.950 ;
        RECT 138.550 192.670 139.450 192.720 ;
        RECT 138.415 192.660 139.450 192.670 ;
        RECT 133.505 191.530 134.565 191.760 ;
        RECT 124.690 189.260 125.460 189.760 ;
        RECT 126.750 189.260 127.550 189.760 ;
        RECT 124.690 188.990 124.920 189.260 ;
        RECT 125.230 188.990 125.460 189.260 ;
        RECT 126.780 188.990 127.010 189.260 ;
        RECT 127.320 188.990 127.550 189.260 ;
        RECT 128.870 188.990 129.150 189.950 ;
        RECT 121.440 188.860 122.440 188.940 ;
        RECT 123.530 188.860 124.530 188.940 ;
        RECT 125.620 188.860 126.620 188.940 ;
        RECT 127.710 188.860 128.710 188.940 ;
        RECT 121.400 188.710 122.440 188.860 ;
        RECT 123.500 188.710 124.530 188.860 ;
        RECT 125.600 188.710 126.620 188.860 ;
        RECT 127.700 188.710 128.710 188.860 ;
        RECT 121.400 188.330 122.400 188.710 ;
        RECT 123.500 188.330 124.500 188.710 ;
        RECT 125.600 188.330 126.600 188.710 ;
        RECT 127.700 188.330 128.700 188.710 ;
        RECT 121.400 188.160 122.440 188.330 ;
        RECT 123.500 188.160 124.530 188.330 ;
        RECT 125.600 188.160 126.620 188.330 ;
        RECT 127.700 188.160 128.710 188.330 ;
        RECT 121.440 188.100 122.440 188.160 ;
        RECT 123.530 188.100 124.530 188.160 ;
        RECT 125.620 188.100 126.620 188.160 ;
        RECT 127.710 188.100 128.710 188.160 ;
        RECT 128.950 188.050 129.150 188.990 ;
        RECT 121.050 187.090 121.280 188.050 ;
        RECT 122.600 187.760 122.830 188.050 ;
        RECT 123.140 187.760 123.370 188.050 ;
        RECT 122.600 187.260 123.370 187.760 ;
        RECT 121.450 187.040 122.350 187.210 ;
        RECT 122.600 187.090 122.830 187.260 ;
        RECT 123.140 187.090 123.370 187.260 ;
        RECT 124.690 187.760 124.920 188.050 ;
        RECT 125.230 187.760 125.460 188.050 ;
        RECT 126.780 187.760 127.010 188.050 ;
        RECT 127.320 187.760 127.550 188.050 ;
        RECT 124.690 187.260 125.460 187.760 ;
        RECT 126.750 187.260 127.550 187.760 ;
        RECT 123.550 187.040 124.450 187.210 ;
        RECT 124.690 187.090 124.920 187.260 ;
        RECT 125.230 187.090 125.460 187.260 ;
        RECT 125.650 187.040 126.550 187.210 ;
        RECT 126.780 187.090 127.010 187.260 ;
        RECT 127.320 187.090 127.550 187.260 ;
        RECT 127.750 187.040 128.650 187.210 ;
        RECT 128.870 187.090 129.150 188.050 ;
        RECT 121.440 186.810 122.440 187.040 ;
        RECT 123.530 186.810 124.530 187.040 ;
        RECT 125.620 186.810 126.620 187.040 ;
        RECT 127.710 186.810 128.710 187.040 ;
        RECT 119.350 185.500 120.580 186.720 ;
        RECT 121.500 186.430 122.400 186.510 ;
        RECT 123.600 186.430 124.500 186.510 ;
        RECT 125.600 186.430 126.600 186.510 ;
        RECT 127.700 186.430 128.700 186.610 ;
        RECT 121.440 186.200 122.440 186.430 ;
        RECT 123.530 186.200 124.530 186.430 ;
        RECT 125.600 186.200 126.620 186.430 ;
        RECT 127.700 186.200 128.710 186.430 ;
        RECT 119.350 182.660 120.400 185.500 ;
        RECT 121.050 185.190 121.280 186.150 ;
        RECT 121.500 186.110 122.400 186.200 ;
        RECT 122.600 185.860 122.830 186.150 ;
        RECT 123.140 185.860 123.370 186.150 ;
        RECT 123.600 186.110 124.500 186.200 ;
        RECT 122.600 185.360 123.370 185.860 ;
        RECT 122.600 185.190 122.830 185.360 ;
        RECT 123.140 185.190 123.370 185.360 ;
        RECT 124.690 185.860 124.920 186.150 ;
        RECT 125.230 185.860 125.460 186.150 ;
        RECT 125.600 186.010 126.600 186.200 ;
        RECT 126.780 185.860 127.010 186.150 ;
        RECT 127.320 185.860 127.550 186.150 ;
        RECT 127.700 186.110 128.700 186.200 ;
        RECT 128.950 186.150 129.150 187.090 ;
        RECT 124.690 185.360 125.460 185.860 ;
        RECT 126.750 185.360 127.550 185.860 ;
        RECT 124.690 185.190 124.920 185.360 ;
        RECT 125.230 185.190 125.460 185.360 ;
        RECT 126.780 185.190 127.010 185.360 ;
        RECT 127.320 185.190 127.550 185.360 ;
        RECT 128.870 185.190 129.150 186.150 ;
        RECT 121.440 184.910 122.440 185.140 ;
        RECT 123.530 184.910 124.530 185.140 ;
        RECT 125.620 184.910 126.620 185.140 ;
        RECT 127.710 184.910 128.710 185.140 ;
        RECT 121.500 184.530 122.400 184.910 ;
        RECT 123.600 184.530 124.500 184.910 ;
        RECT 125.700 184.530 126.600 184.910 ;
        RECT 127.800 184.530 128.700 184.910 ;
        RECT 121.440 184.300 122.440 184.530 ;
        RECT 123.530 184.300 124.530 184.530 ;
        RECT 125.620 184.300 126.620 184.530 ;
        RECT 127.710 184.300 128.710 184.530 ;
        RECT 128.950 184.250 129.150 185.190 ;
        RECT 121.050 183.290 121.280 184.250 ;
        RECT 122.600 184.060 122.830 184.250 ;
        RECT 123.140 184.060 123.370 184.250 ;
        RECT 122.600 183.560 123.370 184.060 ;
        RECT 121.500 183.240 122.400 183.310 ;
        RECT 122.600 183.290 122.830 183.560 ;
        RECT 123.140 183.290 123.370 183.560 ;
        RECT 124.690 184.060 124.920 184.250 ;
        RECT 125.230 184.060 125.460 184.250 ;
        RECT 126.780 184.060 127.010 184.250 ;
        RECT 127.320 184.060 127.550 184.250 ;
        RECT 124.690 183.560 125.460 184.060 ;
        RECT 126.750 183.560 127.550 184.060 ;
        RECT 123.600 183.240 124.500 183.310 ;
        RECT 124.690 183.290 124.920 183.560 ;
        RECT 125.230 183.290 125.460 183.560 ;
        RECT 125.700 183.240 126.600 183.310 ;
        RECT 126.780 183.290 127.010 183.560 ;
        RECT 127.320 183.290 127.550 183.560 ;
        RECT 128.870 183.410 129.150 184.250 ;
        RECT 127.700 183.240 128.600 183.410 ;
        RECT 128.870 183.290 129.250 183.410 ;
        RECT 121.440 183.010 122.440 183.240 ;
        RECT 123.530 183.010 124.530 183.240 ;
        RECT 125.620 183.010 126.620 183.240 ;
        RECT 127.700 183.010 128.710 183.240 ;
        RECT 121.500 182.910 122.400 183.010 ;
        RECT 123.600 182.910 124.500 183.010 ;
        RECT 125.700 182.910 126.600 183.010 ;
        RECT 128.950 182.910 129.250 183.290 ;
        RECT 119.350 182.460 128.850 182.660 ;
        RECT 119.350 182.350 129.050 182.460 ;
        RECT 119.350 181.060 129.100 182.350 ;
        RECT 129.750 181.710 130.150 183.310 ;
        RECT 130.750 183.110 131.150 190.310 ;
        RECT 132.150 190.240 133.795 190.470 ;
        RECT 132.150 187.890 133.350 190.240 ;
        RECT 134.050 189.180 134.550 191.530 ;
        RECT 134.855 190.520 135.085 191.480 ;
        RECT 138.350 190.370 139.450 192.660 ;
        RECT 140.450 191.660 140.850 193.330 ;
        RECT 141.055 191.710 141.285 192.670 ;
        RECT 145.420 192.560 145.680 192.620 ;
        RECT 145.850 192.560 146.850 195.160 ;
        RECT 145.420 191.760 146.850 192.560 ;
        RECT 145.420 191.700 145.680 191.760 ;
        RECT 139.705 191.460 140.850 191.660 ;
        RECT 139.705 191.430 140.765 191.460 ;
        RECT 141.055 190.420 141.285 191.380 ;
        RECT 134.855 189.230 135.085 190.190 ;
        RECT 138.350 190.160 139.995 190.370 ;
        RECT 133.505 188.950 134.565 189.180 ;
        RECT 132.150 187.660 133.795 187.890 ;
        RECT 131.450 181.610 131.750 186.610 ;
        RECT 132.150 185.310 133.350 187.660 ;
        RECT 134.050 186.600 134.550 188.950 ;
        RECT 134.855 187.940 135.085 188.900 ;
        RECT 134.855 186.650 135.085 187.610 ;
        RECT 133.505 186.370 134.565 186.600 ;
        RECT 132.150 185.080 133.795 185.310 ;
        RECT 132.150 182.730 133.350 185.080 ;
        RECT 134.050 184.020 134.550 186.370 ;
        RECT 134.855 185.360 135.085 186.320 ;
        RECT 134.855 184.070 135.085 185.030 ;
        RECT 138.350 184.660 138.650 190.160 ;
        RECT 138.935 190.140 139.995 190.160 ;
        RECT 138.850 189.750 139.350 189.760 ;
        RECT 138.850 189.520 139.995 189.750 ;
        RECT 138.850 187.170 139.350 189.520 ;
        RECT 141.055 188.510 141.285 189.470 ;
        RECT 139.705 188.230 140.850 188.460 ;
        RECT 138.850 186.940 139.995 187.170 ;
        RECT 138.415 184.640 138.645 184.660 ;
        RECT 138.850 184.590 139.350 186.940 ;
        RECT 140.350 185.880 140.850 188.230 ;
        RECT 141.055 187.220 141.285 188.180 ;
        RECT 143.550 187.950 144.150 188.810 ;
        RECT 143.105 187.760 144.165 187.950 ;
        RECT 143.105 187.720 144.650 187.760 ;
        RECT 143.550 187.670 144.650 187.720 ;
        RECT 141.055 185.930 141.285 186.890 ;
        RECT 141.815 186.710 142.045 187.670 ;
        RECT 143.550 187.660 144.685 187.670 ;
        RECT 143.550 186.660 144.750 187.660 ;
        RECT 143.105 186.560 144.750 186.660 ;
        RECT 145.420 186.960 145.680 187.020 ;
        RECT 145.850 186.960 146.850 191.760 ;
        RECT 143.105 186.430 144.165 186.560 ;
        RECT 143.550 186.050 144.150 186.430 ;
        RECT 145.420 186.160 146.850 186.960 ;
        RECT 145.420 186.100 145.680 186.160 ;
        RECT 139.705 185.650 140.850 185.880 ;
        RECT 142.250 185.820 144.250 186.050 ;
        RECT 138.850 184.360 139.995 184.590 ;
        RECT 133.505 183.790 134.565 184.020 ;
        RECT 138.850 183.950 139.350 184.360 ;
        RECT 140.350 184.260 140.850 185.650 ;
        RECT 141.815 185.760 142.045 185.770 ;
        RECT 143.550 185.760 144.150 185.820 ;
        RECT 141.055 184.640 141.285 185.600 ;
        RECT 141.815 184.810 142.050 185.760 ;
        RECT 132.150 182.560 133.795 182.730 ;
        RECT 132.735 182.500 133.795 182.560 ;
        RECT 134.050 182.150 134.550 183.790 ;
        RECT 134.855 182.780 135.085 183.740 ;
        RECT 138.850 183.720 139.995 183.950 ;
        RECT 141.850 183.870 142.050 184.810 ;
        RECT 142.250 184.760 143.350 185.010 ;
        RECT 144.455 184.810 144.685 185.770 ;
        RECT 142.250 184.530 144.250 184.760 ;
        RECT 142.250 184.510 143.350 184.530 ;
        RECT 142.450 184.150 143.150 184.160 ;
        RECT 142.250 183.920 144.250 184.150 ;
        RECT 136.450 183.660 137.050 183.710 ;
        RECT 133.505 181.960 134.565 182.150 ;
        RECT 133.505 181.920 135.150 181.960 ;
        RECT 132.215 180.910 132.445 181.870 ;
        RECT 134.050 180.860 135.150 181.920 ;
        RECT 133.505 180.630 134.565 180.860 ;
        RECT 134.050 180.390 134.550 180.630 ;
        RECT 133.990 179.930 134.610 180.390 ;
        RECT 134.050 176.560 134.550 179.930 ;
        RECT 136.350 176.560 137.050 183.660 ;
        RECT 138.350 183.110 138.650 183.710 ;
        RECT 138.415 182.710 138.650 183.110 ;
        RECT 138.450 182.380 138.650 182.710 ;
        RECT 138.415 181.420 138.650 182.380 ;
        RECT 138.450 181.090 138.650 181.420 ;
        RECT 138.415 180.130 138.650 181.090 ;
        RECT 138.450 179.800 138.650 180.130 ;
        RECT 138.415 178.860 138.650 179.800 ;
        RECT 138.850 181.370 139.350 183.720 ;
        RECT 141.815 183.710 142.050 183.870 ;
        RECT 141.055 182.710 141.285 183.670 ;
        RECT 141.750 183.110 142.050 183.710 ;
        RECT 139.705 182.430 140.765 182.660 ;
        RECT 138.850 181.140 139.995 181.370 ;
        RECT 138.415 178.840 138.645 178.860 ;
        RECT 138.850 178.790 139.350 181.140 ;
        RECT 140.250 180.080 140.750 182.430 ;
        RECT 141.055 181.420 141.285 182.380 ;
        RECT 141.055 180.130 141.285 181.090 ;
        RECT 139.705 179.850 140.765 180.080 ;
        RECT 141.055 178.840 141.285 179.800 ;
        RECT 141.815 178.910 142.045 183.110 ;
        RECT 142.450 179.860 143.150 183.920 ;
        RECT 142.450 179.810 143.050 179.860 ;
        RECT 144.455 178.910 144.685 183.870 ;
        RECT 145.420 183.060 145.680 183.120 ;
        RECT 145.850 183.060 146.850 186.160 ;
        RECT 145.420 182.260 146.850 183.060 ;
        RECT 145.420 182.200 145.680 182.260 ;
        RECT 138.850 178.560 139.995 178.790 ;
        RECT 142.250 178.630 144.250 178.860 ;
        RECT 138.850 178.150 139.350 178.560 ;
        RECT 143.450 178.250 144.150 178.630 ;
        RECT 145.420 178.460 145.680 178.520 ;
        RECT 145.850 178.460 146.850 182.260 ;
        RECT 143.105 178.160 144.165 178.250 ;
        RECT 138.850 177.920 139.995 178.150 ;
        RECT 143.105 178.020 144.550 178.160 ;
        RECT 143.450 177.970 144.550 178.020 ;
        RECT 138.415 177.860 138.645 177.870 ;
        RECT 138.850 177.860 139.350 177.920 ;
        RECT 138.415 176.960 139.350 177.860 ;
        RECT 138.415 176.910 138.645 176.960 ;
        RECT 138.850 176.860 139.350 176.960 ;
        RECT 141.055 176.910 141.285 177.870 ;
        RECT 141.815 177.010 142.045 177.970 ;
        RECT 143.450 177.010 144.685 177.970 ;
        RECT 145.420 177.660 146.850 178.460 ;
        RECT 145.420 177.600 145.680 177.660 ;
        RECT 143.450 176.960 144.650 177.010 ;
        RECT 143.105 176.860 144.650 176.960 ;
        RECT 138.850 176.630 139.995 176.860 ;
        RECT 143.105 176.730 144.165 176.860 ;
        RECT 143.450 176.660 144.150 176.730 ;
        RECT 138.850 176.560 139.350 176.630 ;
        RECT 127.450 169.920 128.450 171.860 ;
        RECT 127.450 168.960 128.460 169.920 ;
        RECT 127.460 168.920 128.460 168.960 ;
        RECT 129.060 168.920 130.060 169.920 ;
        RECT 133.850 168.960 134.850 176.560 ;
        RECT 136.150 174.910 137.150 176.560 ;
        RECT 143.550 176.010 144.150 176.660 ;
        RECT 145.850 175.560 146.850 177.660 ;
        RECT 127.660 156.770 128.260 168.920 ;
        RECT 129.460 161.170 129.860 168.920 ;
        RECT 137.760 167.910 138.660 167.920 ;
        RECT 137.760 167.680 145.675 167.910 ;
        RECT 130.325 167.620 130.555 167.630 ;
        RECT 130.325 166.670 130.560 167.620 ;
        RECT 130.360 166.620 130.560 166.670 ;
        RECT 137.760 166.620 138.660 167.680 ;
        RECT 130.360 166.520 138.660 166.620 ;
        RECT 130.360 166.390 138.405 166.520 ;
        RECT 130.360 166.320 132.060 166.390 ;
        RECT 130.360 164.020 130.560 166.320 ;
        RECT 134.560 164.040 135.060 166.390 ;
        RECT 145.960 166.340 146.160 167.620 ;
        RECT 143.760 165.330 144.960 165.470 ;
        RECT 145.960 165.380 146.195 166.340 ;
        RECT 138.115 165.100 145.675 165.330 ;
        RECT 143.760 164.870 144.960 165.100 ;
        RECT 145.960 165.050 146.160 165.380 ;
        RECT 145.960 164.090 146.195 165.050 ;
        RECT 130.845 164.020 138.405 164.040 ;
        RECT 130.360 163.810 138.660 164.020 ;
        RECT 130.360 163.760 132.060 163.810 ;
        RECT 130.325 163.720 132.060 163.760 ;
        RECT 130.325 162.820 130.560 163.720 ;
        RECT 130.325 162.800 130.555 162.820 ;
        RECT 132.330 155.660 132.790 156.280 ;
        RECT 133.260 152.610 134.060 152.620 ;
        RECT 133.110 151.650 134.060 152.610 ;
        RECT 134.560 152.070 135.060 163.810 ;
        RECT 137.760 162.750 138.660 163.810 ;
        RECT 137.760 162.620 145.675 162.750 ;
        RECT 138.115 162.520 145.675 162.620 ;
        RECT 144.845 162.020 145.405 162.110 ;
        RECT 144.360 161.830 145.560 162.020 ;
        RECT 138.060 158.690 138.460 158.720 ;
        RECT 137.885 158.460 138.460 158.690 ;
        RECT 137.410 158.320 137.640 158.410 ;
        RECT 138.060 158.320 138.460 158.460 ;
        RECT 138.960 158.320 139.190 158.410 ;
        RECT 137.410 157.620 139.190 158.320 ;
        RECT 137.410 157.450 137.640 157.620 ;
        RECT 138.060 157.400 138.460 157.620 ;
        RECT 138.960 157.450 139.190 157.620 ;
        RECT 138.060 157.220 138.715 157.400 ;
        RECT 137.460 157.170 138.715 157.220 ;
        RECT 137.460 157.120 138.460 157.170 ;
        RECT 137.410 156.820 138.460 157.120 ;
        RECT 137.410 156.160 137.660 156.820 ;
        RECT 138.060 156.770 138.460 156.820 ;
        RECT 137.460 155.830 137.660 156.160 ;
        RECT 137.410 154.870 137.660 155.830 ;
        RECT 137.860 156.110 138.360 156.270 ;
        RECT 138.960 156.160 139.190 157.120 ;
        RECT 137.860 155.880 138.445 156.110 ;
        RECT 137.860 155.670 138.360 155.880 ;
        RECT 138.960 154.870 139.190 155.830 ;
        RECT 137.460 154.820 137.660 154.870 ;
        RECT 138.160 154.820 138.660 154.870 ;
        RECT 138.155 154.720 138.715 154.820 ;
        RECT 137.410 154.420 137.640 154.540 ;
        RECT 138.060 154.420 138.760 154.720 ;
        RECT 138.960 154.420 139.190 154.540 ;
        RECT 137.410 153.580 139.190 154.420 ;
        RECT 137.460 153.420 139.160 153.580 ;
        RECT 137.885 153.300 138.445 153.420 ;
        RECT 135.560 152.890 136.160 152.920 ;
        RECT 135.560 152.820 138.415 152.890 ;
        RECT 135.560 152.660 138.860 152.820 ;
        RECT 133.260 151.600 134.060 151.650 ;
        RECT 135.560 151.600 136.160 152.660 ;
        RECT 138.160 152.610 138.860 152.660 ;
        RECT 133.260 151.520 136.160 151.600 ;
        RECT 133.585 151.420 136.160 151.520 ;
        RECT 133.585 151.370 136.145 151.420 ;
        RECT 133.110 150.360 133.340 151.320 ;
        RECT 132.330 148.560 132.790 149.180 ;
        RECT 133.110 149.070 133.340 150.030 ;
        RECT 134.460 149.170 134.960 151.370 ;
        RECT 137.360 151.220 137.860 152.520 ;
        RECT 138.160 151.720 138.890 152.610 ;
        RECT 139.360 152.370 139.660 154.870 ;
        RECT 138.660 151.650 138.890 151.720 ;
        RECT 138.660 151.220 138.890 151.320 ;
        RECT 137.360 150.310 138.960 151.220 ;
        RECT 139.860 150.820 140.160 161.570 ;
        RECT 144.325 160.870 145.560 161.830 ;
        RECT 144.360 160.820 145.560 160.870 ;
        RECT 144.360 160.720 145.760 160.820 ;
        RECT 145.115 160.590 145.760 160.720 ;
        RECT 144.325 160.520 144.555 160.540 ;
        RECT 144.325 159.580 144.560 160.520 ;
        RECT 144.360 159.250 144.560 159.580 ;
        RECT 144.325 158.290 144.560 159.250 ;
        RECT 144.360 157.960 144.560 158.290 ;
        RECT 144.325 157.000 144.560 157.960 ;
        RECT 144.360 156.670 144.560 157.000 ;
        RECT 144.325 155.710 144.560 156.670 ;
        RECT 144.360 155.420 144.560 155.710 ;
        RECT 144.760 159.530 144.960 159.620 ;
        RECT 144.760 159.300 145.405 159.530 ;
        RECT 144.760 156.950 144.960 159.300 ;
        RECT 145.560 158.240 145.760 160.590 ;
        RECT 145.960 160.540 146.160 164.090 ;
        RECT 145.960 159.620 146.195 160.540 ;
        RECT 145.965 159.580 146.195 159.620 ;
        RECT 145.115 158.010 145.760 158.240 ;
        RECT 144.760 156.720 145.405 156.950 ;
        RECT 144.760 155.420 144.960 156.720 ;
        RECT 145.560 155.870 145.760 158.010 ;
        RECT 145.360 155.660 145.760 155.870 ;
        RECT 145.115 155.430 145.760 155.660 ;
        RECT 144.360 155.380 144.960 155.420 ;
        RECT 144.325 154.470 144.960 155.380 ;
        RECT 145.360 155.270 145.760 155.430 ;
        RECT 141.960 153.620 142.360 154.470 ;
        RECT 144.325 154.420 145.260 154.470 ;
        RECT 144.760 154.370 145.260 154.420 ;
        RECT 146.460 154.420 147.160 165.420 ;
        RECT 153.650 162.060 155.350 162.260 ;
        RECT 153.650 160.460 157.050 162.060 ;
        RECT 153.650 160.260 155.350 160.460 ;
        RECT 144.760 154.220 145.405 154.370 ;
        RECT 144.360 154.090 145.760 154.220 ;
        RECT 140.960 153.420 142.360 153.620 ;
        RECT 140.460 153.020 142.360 153.420 ;
        RECT 144.325 153.130 145.760 154.090 ;
        RECT 141.505 152.880 142.315 153.020 ;
        RECT 140.960 152.630 141.360 152.770 ;
        RECT 140.460 152.120 140.760 152.420 ;
        RECT 140.960 152.400 141.795 152.630 ;
        RECT 142.560 152.470 142.860 152.970 ;
        RECT 140.960 152.370 141.360 152.400 ;
        RECT 140.460 151.270 140.660 152.120 ;
        RECT 141.505 152.020 142.315 152.150 ;
        RECT 141.260 151.940 142.660 152.020 ;
        RECT 141.260 151.920 142.790 151.940 ;
        RECT 141.260 151.670 142.860 151.920 ;
        RECT 140.985 151.620 142.860 151.670 ;
        RECT 140.985 151.520 142.660 151.620 ;
        RECT 140.985 151.440 141.795 151.520 ;
        RECT 140.460 150.870 140.760 151.270 ;
        RECT 140.460 150.820 140.660 150.870 ;
        RECT 141.960 150.770 142.360 151.520 ;
        RECT 135.855 150.220 138.960 150.310 ;
        RECT 135.855 150.080 138.415 150.220 ;
        RECT 133.660 149.020 134.960 149.170 ;
        RECT 133.585 148.790 136.145 149.020 ;
        RECT 133.660 148.770 134.960 148.790 ;
        RECT 133.110 147.780 133.340 148.740 ;
        RECT 133.110 146.490 133.340 147.450 ;
        RECT 134.460 146.440 134.960 148.770 ;
        RECT 135.855 147.500 138.415 147.730 ;
        RECT 133.585 146.420 136.145 146.440 ;
        RECT 133.585 146.320 136.160 146.420 ;
        RECT 133.160 146.210 136.160 146.320 ;
        RECT 133.160 146.160 133.860 146.210 ;
        RECT 133.110 145.420 133.860 146.160 ;
        RECT 134.960 145.720 135.260 145.770 ;
        RECT 133.110 145.200 133.340 145.420 ;
        RECT 130.360 142.630 130.660 142.720 ;
        RECT 130.325 141.670 130.660 142.630 ;
        RECT 130.360 141.620 130.660 141.670 ;
        RECT 134.960 141.620 135.360 145.720 ;
        RECT 135.860 145.150 136.160 146.210 ;
        RECT 136.760 145.420 137.260 147.500 ;
        RECT 138.660 146.520 138.960 150.220 ;
        RECT 138.660 146.490 138.890 146.520 ;
        RECT 138.660 146.120 138.890 146.160 ;
        RECT 137.960 145.200 138.890 146.120 ;
        RECT 137.960 145.150 138.860 145.200 ;
        RECT 135.855 145.020 138.860 145.150 ;
        RECT 135.855 144.920 138.415 145.020 ;
        RECT 143.060 143.670 143.460 152.970 ;
        RECT 144.360 152.920 145.760 153.130 ;
        RECT 146.460 153.020 147.060 154.420 ;
        RECT 146.460 153.010 148.060 153.020 ;
        RECT 145.115 152.850 145.675 152.920 ;
        RECT 144.845 152.320 145.405 152.510 ;
        RECT 144.360 152.130 145.560 152.320 ;
        RECT 144.325 151.220 145.560 152.130 ;
        RECT 146.460 151.910 148.850 153.010 ;
        RECT 144.325 151.170 145.675 151.220 ;
        RECT 144.360 151.120 145.675 151.170 ;
        RECT 144.360 151.020 145.760 151.120 ;
        RECT 144.360 150.840 144.860 151.020 ;
        RECT 145.115 150.990 145.760 151.020 ;
        RECT 144.325 150.720 144.860 150.840 ;
        RECT 145.160 150.770 145.760 150.990 ;
        RECT 144.325 149.880 144.560 150.720 ;
        RECT 144.360 149.550 144.560 149.880 ;
        RECT 144.325 148.590 144.560 149.550 ;
        RECT 144.360 148.260 144.560 148.590 ;
        RECT 144.325 147.300 144.560 148.260 ;
        RECT 144.360 146.970 144.560 147.300 ;
        RECT 144.325 146.010 144.560 146.970 ;
        RECT 144.360 145.780 144.560 146.010 ;
        RECT 144.325 144.920 144.560 145.780 ;
        RECT 144.760 149.930 145.360 150.070 ;
        RECT 144.760 149.700 145.405 149.930 ;
        RECT 144.760 149.570 145.360 149.700 ;
        RECT 144.760 147.350 144.960 149.570 ;
        RECT 145.560 148.640 145.760 150.770 ;
        RECT 145.115 148.410 145.760 148.640 ;
        RECT 144.760 147.120 145.405 147.350 ;
        RECT 144.325 144.820 144.555 144.920 ;
        RECT 144.760 144.770 144.960 147.120 ;
        RECT 145.560 146.060 145.760 148.410 ;
        RECT 145.115 145.830 145.760 146.060 ;
        RECT 145.560 145.820 145.760 145.830 ;
        RECT 144.760 144.540 145.405 144.770 ;
        RECT 144.760 144.520 145.360 144.540 ;
        RECT 144.460 144.490 145.360 144.520 ;
        RECT 144.325 144.020 145.360 144.490 ;
        RECT 144.325 143.480 145.660 144.020 ;
        RECT 144.325 143.430 145.675 143.480 ;
        RECT 144.360 143.320 145.675 143.430 ;
        RECT 145.115 143.250 145.675 143.320 ;
        RECT 145.160 143.220 145.660 143.250 ;
        RECT 137.660 142.910 138.560 142.920 ;
        RECT 137.660 142.680 145.675 142.910 ;
        RECT 137.660 141.620 138.560 142.680 ;
        RECT 130.360 141.420 138.560 141.620 ;
        RECT 130.360 141.390 138.405 141.420 ;
        RECT 130.360 141.320 131.660 141.390 ;
        RECT 130.360 139.020 130.660 141.320 ;
        RECT 134.960 139.040 135.360 141.390 ;
        RECT 142.760 140.330 145.560 140.470 ;
        RECT 138.115 140.100 145.675 140.330 ;
        RECT 142.760 140.070 145.560 140.100 ;
        RECT 137.660 139.040 138.560 139.120 ;
        RECT 130.845 139.020 138.560 139.040 ;
        RECT 130.360 138.810 138.560 139.020 ;
        RECT 130.360 138.760 131.660 138.810 ;
        RECT 130.325 138.720 131.660 138.760 ;
        RECT 130.325 137.820 130.660 138.720 ;
        RECT 130.325 137.800 130.555 137.820 ;
        RECT 134.960 136.620 135.360 138.810 ;
        RECT 137.660 137.750 138.560 138.810 ;
        RECT 145.960 137.820 146.260 145.820 ;
        RECT 146.460 139.920 147.060 151.910 ;
        RECT 137.660 137.620 145.675 137.750 ;
        RECT 138.115 137.520 145.675 137.620 ;
        RECT 134.660 135.620 135.660 136.620 ;
        RECT 123.950 131.360 124.850 131.410 ;
        RECT 121.150 124.260 122.150 125.260 ;
        RECT 123.950 124.260 124.950 131.360 ;
        RECT 127.250 125.260 128.250 126.830 ;
        RECT 125.650 124.660 126.650 125.260 ;
        RECT 125.450 124.260 126.650 124.660 ;
        RECT 127.150 124.260 128.250 125.260 ;
        RECT 140.050 124.260 141.050 125.260 ;
        RECT 145.450 124.360 146.450 136.660 ;
        RECT 119.350 118.160 120.150 123.860 ;
        RECT 121.550 119.710 121.850 124.260 ;
        RECT 119.350 117.160 120.350 118.160 ;
        RECT 119.350 116.610 120.150 117.160 ;
        RECT 119.250 115.810 120.150 116.610 ;
        RECT 119.350 109.660 120.150 115.810 ;
        RECT 122.650 111.510 122.950 122.310 ;
        RECT 123.150 113.190 123.630 123.770 ;
        RECT 124.450 123.690 124.750 124.260 ;
        RECT 125.450 124.160 126.350 124.260 ;
        RECT 124.390 123.430 124.810 123.690 ;
        RECT 125.850 123.560 126.350 124.160 ;
        RECT 124.465 122.930 124.695 123.220 ;
        RECT 124.000 121.860 124.350 122.360 ;
        RECT 124.510 121.385 124.650 122.930 ;
        RECT 125.145 122.525 125.375 122.815 ;
        RECT 124.465 121.095 124.695 121.385 ;
        RECT 124.050 120.025 124.350 120.110 ;
        RECT 124.050 119.710 124.355 120.025 ;
        RECT 124.125 119.375 124.355 119.710 ;
        RECT 124.170 116.725 124.310 119.375 ;
        RECT 124.510 117.805 124.650 121.095 ;
        RECT 125.190 120.925 125.330 122.525 ;
        RECT 125.145 120.635 125.375 120.925 ;
        RECT 125.190 117.805 125.330 120.635 ;
        RECT 124.465 117.515 124.695 117.805 ;
        RECT 125.145 117.515 125.375 117.805 ;
        RECT 124.170 116.435 124.670 116.725 ;
        RECT 124.170 116.425 124.355 116.435 ;
        RECT 124.125 116.135 124.355 116.425 ;
        RECT 123.820 114.700 124.180 115.120 ;
        RECT 123.850 112.410 124.150 114.700 ;
        RECT 124.420 113.250 124.680 113.570 ;
        RECT 124.450 112.310 124.650 113.250 ;
        RECT 125.870 113.190 126.350 123.560 ;
        RECT 124.350 111.810 124.750 112.310 ;
        RECT 127.350 111.860 127.900 124.260 ;
        RECT 139.350 123.960 141.450 124.260 ;
        RECT 146.050 123.960 148.050 124.060 ;
        RECT 135.250 123.710 137.250 123.810 ;
        RECT 130.980 123.460 133.085 123.710 ;
        RECT 135.135 123.460 137.250 123.710 ;
        RECT 131.050 122.880 132.950 123.460 ;
        RECT 135.250 123.410 137.250 123.460 ;
        RECT 130.980 122.630 133.085 122.880 ;
        RECT 135.135 122.630 137.240 122.880 ;
        RECT 135.250 122.050 137.150 122.630 ;
        RECT 130.980 121.800 133.085 122.050 ;
        RECT 135.135 121.800 137.240 122.050 ;
        RECT 131.050 121.220 132.950 121.800 ;
        RECT 130.980 120.970 133.085 121.220 ;
        RECT 135.135 120.970 137.240 121.220 ;
        RECT 135.250 120.390 137.150 120.970 ;
        RECT 130.980 120.140 133.085 120.390 ;
        RECT 135.135 120.140 137.240 120.390 ;
        RECT 131.050 119.560 132.950 120.140 ;
        RECT 130.980 119.310 133.085 119.560 ;
        RECT 135.135 119.310 137.240 119.560 ;
        RECT 135.250 118.730 137.150 119.310 ;
        RECT 130.980 118.480 133.085 118.730 ;
        RECT 135.135 118.480 137.240 118.730 ;
        RECT 131.050 117.900 132.950 118.480 ;
        RECT 130.980 117.650 133.085 117.900 ;
        RECT 135.135 117.650 137.240 117.900 ;
        RECT 132.050 114.560 132.550 114.610 ;
        RECT 122.600 111.410 122.950 111.510 ;
        RECT 121.750 111.110 122.950 111.410 ;
        RECT 121.750 110.970 122.650 111.110 ;
        RECT 125.250 110.970 128.150 111.410 ;
        RECT 121.350 110.780 121.550 110.860 ;
        RECT 121.330 110.490 121.560 110.780 ;
        RECT 121.720 110.740 122.720 110.970 ;
        RECT 125.115 110.860 128.150 110.970 ;
        RECT 122.950 110.810 123.150 110.860 ;
        RECT 124.650 110.810 124.850 110.860 ;
        RECT 122.950 110.780 123.250 110.810 ;
        RECT 121.350 110.460 121.550 110.490 ;
        RECT 121.720 110.300 122.720 110.530 ;
        RECT 122.880 110.490 123.250 110.780 ;
        RECT 122.950 110.410 123.250 110.490 ;
        RECT 124.550 110.780 124.850 110.810 ;
        RECT 124.550 110.490 124.910 110.780 ;
        RECT 125.115 110.740 128.115 110.860 ;
        RECT 128.350 110.780 128.650 110.910 ;
        RECT 124.550 110.410 124.850 110.490 ;
        RECT 125.115 110.300 128.115 110.530 ;
        RECT 128.320 110.510 128.650 110.780 ;
        RECT 128.320 110.490 128.550 110.510 ;
        RECT 128.350 110.460 128.550 110.490 ;
        RECT 121.750 110.060 122.650 110.300 ;
        RECT 119.450 109.610 120.050 109.660 ;
        RECT 121.650 109.460 122.650 110.060 ;
        RECT 125.250 109.990 128.050 110.300 ;
        RECT 125.190 109.730 128.110 109.990 ;
        RECT 125.250 109.560 128.050 109.730 ;
        RECT 125.550 109.510 125.950 109.560 ;
        RECT 126.250 109.510 126.650 109.560 ;
        RECT 126.950 109.510 127.350 109.560 ;
        RECT 127.550 109.510 127.950 109.560 ;
        RECT 131.950 77.960 132.550 114.560 ;
        RECT 135.450 114.060 136.650 117.650 ;
        RECT 135.450 114.010 136.550 114.060 ;
        RECT 137.850 110.910 138.350 123.910 ;
        RECT 139.320 123.710 141.450 123.960 ;
        RECT 145.975 123.710 148.080 123.960 ;
        RECT 139.350 123.660 141.450 123.710 ;
        RECT 139.350 123.130 141.350 123.160 ;
        RECT 146.050 123.130 148.050 123.710 ;
        RECT 139.320 122.880 141.425 123.130 ;
        RECT 145.975 122.880 148.080 123.130 ;
        RECT 139.350 122.300 141.350 122.880 ;
        RECT 139.320 122.050 141.425 122.300 ;
        RECT 145.975 122.050 148.080 122.300 ;
        RECT 146.050 121.470 148.050 122.050 ;
        RECT 139.320 121.220 141.425 121.470 ;
        RECT 145.975 121.220 148.080 121.470 ;
        RECT 139.350 120.640 141.350 121.220 ;
        RECT 146.050 121.160 148.050 121.220 ;
        RECT 146.050 120.640 148.050 120.660 ;
        RECT 139.320 120.390 141.425 120.640 ;
        RECT 145.975 120.390 148.080 120.640 ;
        RECT 139.350 120.360 141.350 120.390 ;
        RECT 139.350 119.810 141.350 119.860 ;
        RECT 146.050 119.810 148.050 120.390 ;
        RECT 139.320 119.560 141.425 119.810 ;
        RECT 145.975 119.560 148.080 119.810 ;
        RECT 139.350 118.980 141.350 119.560 ;
        RECT 139.320 118.730 141.425 118.980 ;
        RECT 145.975 118.730 148.080 118.980 ;
        RECT 146.050 118.150 148.050 118.730 ;
        RECT 139.320 117.900 141.425 118.150 ;
        RECT 145.975 117.900 148.080 118.150 ;
        RECT 139.350 116.590 141.350 117.900 ;
        RECT 146.050 117.860 148.050 117.900 ;
        RECT 139.320 116.340 141.425 116.590 ;
        RECT 145.975 116.340 148.080 116.590 ;
        RECT 146.050 115.760 148.050 116.340 ;
        RECT 139.320 115.510 141.425 115.760 ;
        RECT 145.975 115.510 148.080 115.760 ;
        RECT 139.350 114.930 141.350 115.510 ;
        RECT 146.050 115.460 148.050 115.510 ;
        RECT 139.320 114.680 141.425 114.930 ;
        RECT 145.975 114.680 148.080 114.930 ;
        RECT 139.350 114.560 141.350 114.680 ;
        RECT 146.050 114.100 148.050 114.680 ;
        RECT 139.320 113.850 141.425 114.100 ;
        RECT 145.975 113.850 148.080 114.100 ;
        RECT 139.350 113.270 141.350 113.850 ;
        RECT 146.050 113.760 148.050 113.850 ;
        RECT 139.320 113.020 141.425 113.270 ;
        RECT 145.975 113.020 148.080 113.270 ;
        RECT 139.350 112.960 141.350 113.020 ;
        RECT 137.850 110.210 138.450 110.910 ;
        RECT 138.750 110.860 139.150 112.960 ;
        RECT 139.350 112.440 141.350 112.460 ;
        RECT 146.050 112.440 148.050 113.020 ;
        RECT 139.320 112.190 141.425 112.440 ;
        RECT 145.975 112.190 148.080 112.440 ;
        RECT 139.350 111.610 141.350 112.190 ;
        RECT 146.050 112.160 148.050 112.190 ;
        RECT 139.320 111.360 141.425 111.610 ;
        RECT 145.975 111.360 148.080 111.610 ;
        RECT 138.750 110.780 139.550 110.860 ;
        RECT 146.050 110.780 148.050 111.360 ;
        RECT 138.750 110.530 141.425 110.780 ;
        RECT 145.975 110.530 148.080 110.780 ;
        RECT 138.750 110.460 139.550 110.530 ;
        RECT 146.050 110.460 148.050 110.530 ;
        RECT 147.850 110.060 148.750 110.210 ;
        RECT 146.550 109.460 148.750 110.060 ;
        RECT 146.550 109.410 146.950 109.460 ;
        RECT 147.750 109.060 148.750 109.460 ;
        RECT 131.750 76.860 132.850 77.960 ;
        RECT 131.950 74.610 132.550 76.860 ;
      LAYER via ;
        RECT 109.770 194.470 111.270 195.770 ;
        RECT 107.870 173.970 108.370 174.970 ;
        RECT 107.850 170.960 108.550 171.960 ;
        RECT 119.550 194.360 120.150 195.760 ;
        RECT 121.500 193.760 122.400 194.060 ;
        RECT 123.600 193.760 124.500 194.060 ;
        RECT 125.600 193.760 126.600 194.060 ;
        RECT 127.800 193.760 128.700 194.060 ;
        RECT 130.550 193.760 130.950 194.060 ;
        RECT 119.800 192.060 120.300 192.560 ;
        RECT 121.500 191.960 122.400 192.660 ;
        RECT 123.500 191.960 124.500 192.660 ;
        RECT 125.600 191.960 126.600 192.660 ;
        RECT 127.700 191.960 128.700 192.660 ;
        RECT 121.500 190.560 122.400 190.860 ;
        RECT 123.600 190.560 124.500 190.860 ;
        RECT 125.700 190.560 126.600 190.860 ;
        RECT 127.800 190.560 128.700 190.860 ;
        RECT 121.500 189.960 122.300 190.260 ;
        RECT 123.600 189.960 124.400 190.260 ;
        RECT 125.700 189.960 126.500 190.260 ;
        RECT 127.800 189.960 128.600 190.260 ;
        RECT 140.450 194.760 140.850 195.160 ;
        RECT 145.850 194.760 146.350 195.160 ;
        RECT 130.550 192.060 130.850 192.560 ;
        RECT 130.550 190.560 130.950 190.860 ;
        RECT 138.350 192.060 138.650 192.560 ;
        RECT 119.700 188.260 120.400 188.860 ;
        RECT 121.500 188.260 122.200 188.760 ;
        RECT 123.600 188.260 124.300 188.760 ;
        RECT 125.700 188.260 126.400 188.760 ;
        RECT 127.800 188.360 128.500 188.860 ;
        RECT 121.450 186.860 122.350 187.160 ;
        RECT 123.550 186.860 124.450 187.160 ;
        RECT 125.650 186.860 126.550 187.160 ;
        RECT 127.750 186.860 128.650 187.160 ;
        RECT 121.500 186.160 122.400 186.460 ;
        RECT 123.600 186.160 124.500 186.460 ;
        RECT 125.600 186.060 126.600 186.460 ;
        RECT 127.700 186.160 128.700 186.560 ;
        RECT 119.700 184.360 120.400 185.060 ;
        RECT 121.500 184.460 122.300 185.060 ;
        RECT 123.600 184.460 124.400 185.060 ;
        RECT 125.700 184.460 126.500 185.060 ;
        RECT 127.800 184.460 128.600 185.060 ;
        RECT 121.500 182.960 122.400 183.260 ;
        RECT 123.600 182.960 124.500 183.260 ;
        RECT 130.750 189.960 131.150 190.260 ;
        RECT 130.750 186.760 131.150 187.060 ;
        RECT 125.700 182.960 126.600 183.260 ;
        RECT 127.700 183.060 128.600 183.360 ;
        RECT 128.950 182.960 129.250 183.360 ;
        RECT 129.750 182.960 130.150 183.260 ;
        RECT 130.750 183.160 131.150 183.660 ;
        RECT 131.450 186.260 131.750 186.560 ;
        RECT 129.750 181.760 130.150 182.160 ;
        RECT 143.550 188.160 144.150 188.760 ;
        RECT 145.850 188.160 146.350 188.760 ;
        RECT 140.350 184.560 140.850 184.960 ;
        RECT 132.250 183.260 133.250 183.660 ;
        RECT 131.450 181.660 131.750 182.160 ;
        RECT 142.250 184.560 143.350 184.960 ;
        RECT 136.450 183.160 137.050 183.660 ;
        RECT 134.050 179.760 134.550 180.360 ;
        RECT 138.350 183.160 138.650 183.660 ;
        RECT 141.750 183.160 142.050 183.660 ;
        RECT 140.250 181.660 140.750 182.160 ;
        RECT 145.950 176.760 146.750 179.260 ;
        RECT 143.550 176.060 144.150 176.560 ;
        RECT 145.850 176.060 146.350 176.560 ;
        RECT 133.850 173.960 134.850 174.860 ;
        RECT 127.550 171.160 128.350 171.760 ;
        RECT 129.150 169.060 129.950 169.860 ;
        RECT 133.950 169.060 134.750 169.860 ;
        RECT 143.760 164.920 144.960 165.420 ;
        RECT 146.560 165.020 147.160 165.320 ;
        RECT 129.460 161.220 129.860 161.520 ;
        RECT 127.660 156.820 128.260 157.220 ;
        RECT 110.760 155.820 111.060 156.120 ;
        RECT 132.360 155.720 132.760 156.220 ;
        RECT 139.860 161.220 140.160 161.520 ;
        RECT 138.060 156.820 138.460 157.220 ;
        RECT 137.860 155.720 138.360 156.220 ;
        RECT 138.160 154.520 138.660 154.820 ;
        RECT 139.360 154.420 139.660 154.820 ;
        RECT 134.660 152.120 134.960 152.420 ;
        RECT 137.460 152.120 137.760 152.420 ;
        RECT 110.760 148.720 111.060 149.020 ;
        RECT 107.970 130.470 108.470 131.270 ;
        RECT 107.970 127.570 108.370 128.170 ;
        RECT 107.870 125.870 108.470 126.670 ;
        RECT 107.970 124.370 108.470 125.170 ;
        RECT 132.360 148.620 132.760 149.120 ;
        RECT 139.360 152.420 139.660 152.720 ;
        RECT 145.360 155.320 145.760 155.820 ;
        RECT 153.750 160.460 155.150 162.060 ;
        RECT 146.560 155.320 147.060 155.820 ;
        RECT 141.960 154.020 142.360 154.420 ;
        RECT 144.760 154.020 145.260 154.420 ;
        RECT 140.960 152.420 141.360 152.720 ;
        RECT 142.560 152.520 142.860 152.920 ;
        RECT 143.060 152.520 143.460 152.920 ;
        RECT 137.460 150.720 138.360 151.020 ;
        RECT 139.860 150.920 140.160 151.220 ;
        RECT 140.460 150.920 140.760 151.220 ;
        RECT 141.960 150.820 142.360 151.220 ;
        RECT 133.660 148.820 134.860 149.120 ;
        RECT 134.960 145.420 135.260 145.720 ;
        RECT 136.860 145.520 137.160 145.820 ;
        RECT 135.060 143.820 135.360 144.120 ;
        RECT 147.050 151.960 148.850 152.960 ;
        RECT 145.160 150.820 145.560 151.220 ;
        RECT 144.760 149.620 145.360 150.020 ;
        RECT 146.560 149.620 147.060 150.120 ;
        RECT 143.060 143.720 143.460 144.120 ;
        RECT 142.760 140.120 145.560 140.420 ;
        RECT 146.460 140.120 146.960 140.420 ;
        RECT 134.750 135.760 135.550 136.560 ;
        RECT 145.550 135.760 146.350 136.560 ;
        RECT 123.950 130.460 124.850 131.360 ;
        RECT 121.150 124.460 122.050 125.060 ;
        RECT 145.550 127.560 146.350 128.160 ;
        RECT 127.250 125.960 128.250 126.660 ;
        RECT 125.750 124.460 126.450 125.060 ;
        RECT 140.150 124.460 140.950 125.160 ;
        RECT 145.550 124.560 146.350 125.260 ;
        RECT 109.970 117.370 111.170 118.370 ;
        RECT 119.450 123.260 120.150 123.760 ;
        RECT 123.150 123.260 123.550 123.660 ;
        RECT 121.550 119.760 121.850 120.060 ;
        RECT 122.650 121.960 122.950 122.260 ;
        RECT 119.450 117.260 120.050 118.560 ;
        RECT 124.000 121.910 124.350 122.310 ;
        RECT 124.050 119.760 124.350 120.060 ;
        RECT 123.850 112.460 124.150 112.860 ;
        RECT 124.350 111.860 124.750 112.260 ;
        RECT 135.250 123.460 137.250 123.760 ;
        RECT 137.850 123.360 138.350 123.860 ;
        RECT 127.350 111.910 127.900 112.260 ;
        RECT 132.050 113.960 132.550 114.560 ;
        RECT 137.950 117.060 138.350 117.460 ;
        RECT 122.600 111.160 122.900 111.460 ;
        RECT 125.250 111.060 128.150 111.360 ;
        RECT 122.950 110.460 123.250 110.760 ;
        RECT 124.550 110.460 124.850 110.760 ;
        RECT 128.350 110.560 128.650 110.860 ;
        RECT 131.950 110.460 132.550 110.860 ;
        RECT 119.450 109.660 120.050 110.160 ;
        RECT 121.750 109.660 122.450 110.160 ;
        RECT 125.550 109.560 125.950 109.960 ;
        RECT 126.250 109.560 126.650 109.960 ;
        RECT 126.950 109.560 127.350 109.960 ;
        RECT 127.550 109.560 127.950 109.960 ;
        RECT 139.450 117.060 141.250 117.460 ;
        RECT 138.750 112.460 139.050 112.860 ;
        RECT 137.850 110.260 138.450 110.860 ;
        RECT 147.850 109.260 148.750 110.160 ;
        RECT 131.850 76.960 132.750 77.860 ;
      LAYER met2 ;
        RECT 49.100 196.200 50.500 196.250 ;
        RECT 49.100 195.960 112.700 196.200 ;
        RECT 49.100 194.400 120.250 195.960 ;
        RECT 140.400 194.760 146.400 195.160 ;
        RECT 109.570 194.270 120.250 194.400 ;
        RECT 110.680 194.260 120.250 194.270 ;
        RECT 121.400 193.760 131.000 194.060 ;
        RECT 119.700 191.960 128.750 192.660 ;
        RECT 130.500 192.060 138.700 192.560 ;
        RECT 121.400 190.560 131.000 190.860 ;
        RECT 121.400 189.960 131.200 190.260 ;
        RECT 119.650 188.260 128.600 188.860 ;
        RECT 143.500 188.160 146.400 188.760 ;
        RECT 121.400 187.060 122.400 187.160 ;
        RECT 123.500 187.060 124.500 187.160 ;
        RECT 125.600 187.060 126.600 187.160 ;
        RECT 127.700 187.060 128.700 187.160 ;
        RECT 121.400 186.760 131.200 187.060 ;
        RECT 121.100 186.260 131.800 186.560 ;
        RECT 121.450 186.160 122.450 186.260 ;
        RECT 123.550 186.160 124.550 186.260 ;
        RECT 125.550 186.060 126.650 186.260 ;
        RECT 127.650 186.160 128.750 186.260 ;
        RECT 119.650 184.360 128.700 185.060 ;
        RECT 140.300 184.560 143.400 184.960 ;
        RECT 127.650 183.260 128.650 183.360 ;
        RECT 128.900 183.260 129.300 183.360 ;
        RECT 121.200 182.960 130.200 183.260 ;
        RECT 130.700 183.160 142.100 183.660 ;
        RECT 129.700 181.760 140.800 182.160 ;
        RECT 131.300 181.660 140.800 181.760 ;
        RECT 134.000 179.760 143.150 180.360 ;
        RECT 145.900 176.760 146.800 179.260 ;
        RECT 143.500 176.060 146.400 176.560 ;
        RECT 90.250 174.970 108.800 175.000 ;
        RECT 90.250 174.960 112.430 174.970 ;
        RECT 90.250 173.970 135.020 174.960 ;
        RECT 90.250 173.900 108.800 173.970 ;
        RECT 111.180 173.960 135.020 173.970 ;
        RECT 96.400 171.860 108.600 172.000 ;
        RECT 96.400 171.060 128.450 171.860 ;
        RECT 96.400 171.000 108.600 171.060 ;
        RECT 107.800 170.960 108.600 171.000 ;
        RECT 129.050 168.960 134.850 169.960 ;
        RECT 143.710 165.320 147.160 165.420 ;
        RECT 143.710 165.020 147.210 165.320 ;
        RECT 143.710 164.920 147.160 165.020 ;
        RECT 129.410 161.220 140.210 161.520 ;
        RECT 153.700 160.460 155.200 162.060 ;
        RECT 127.610 156.820 138.510 157.220 ;
        RECT 110.660 155.720 138.410 156.220 ;
        RECT 145.310 155.320 147.110 155.820 ;
        RECT 138.110 154.520 139.710 154.820 ;
        RECT 138.160 154.420 139.710 154.520 ;
        RECT 141.910 154.020 145.360 154.420 ;
        RECT 134.560 152.020 137.860 152.520 ;
        RECT 139.310 152.420 141.410 152.720 ;
        RECT 142.510 152.520 143.510 152.920 ;
        RECT 147.000 151.960 148.900 152.960 ;
        RECT 129.210 151.120 130.710 151.720 ;
        RECT 129.210 151.020 138.360 151.120 ;
        RECT 129.210 150.720 138.410 151.020 ;
        RECT 139.760 150.920 140.810 151.220 ;
        RECT 139.760 150.820 140.660 150.920 ;
        RECT 141.910 150.820 145.610 151.220 ;
        RECT 129.210 150.620 138.360 150.720 ;
        RECT 129.210 149.620 130.710 150.620 ;
        RECT 144.760 150.020 147.110 150.120 ;
        RECT 144.710 149.620 147.110 150.020 ;
        RECT 110.660 148.620 134.960 149.120 ;
        RECT 134.960 145.720 137.210 145.820 ;
        RECT 134.910 145.520 137.210 145.720 ;
        RECT 134.910 145.420 137.160 145.520 ;
        RECT 128.260 144.120 129.760 145.120 ;
        RECT 128.260 143.720 143.510 144.120 ;
        RECT 128.260 142.720 129.760 143.720 ;
        RECT 142.560 140.020 147.060 140.520 ;
        RECT 134.650 135.660 146.450 136.660 ;
        RECT 103.200 131.370 108.400 131.400 ;
        RECT 103.200 131.360 112.430 131.370 ;
        RECT 103.200 130.400 124.950 131.360 ;
        RECT 107.870 130.370 124.950 130.400 ;
        RECT 111.250 130.360 124.950 130.370 ;
        RECT 103.200 128.270 108.900 128.400 ;
        RECT 103.200 128.260 112.430 128.270 ;
        RECT 103.200 127.470 146.450 128.260 ;
        RECT 103.200 127.400 108.900 127.470 ;
        RECT 111.250 127.460 146.450 127.470 ;
        RECT 88.000 126.670 108.000 126.700 ;
        RECT 88.000 126.660 112.430 126.670 ;
        RECT 88.000 125.960 128.300 126.660 ;
        RECT 88.000 125.870 128.250 125.960 ;
        RECT 88.000 125.700 108.000 125.870 ;
        RECT 111.250 125.860 128.250 125.870 ;
        RECT 1.000 125.400 2.400 125.450 ;
        RECT 0.950 125.270 108.150 125.400 ;
        RECT 0.950 125.260 112.430 125.270 ;
        RECT 0.950 124.300 126.650 125.260 ;
        RECT 140.050 124.460 146.450 125.360 ;
        RECT 1.000 124.250 2.400 124.300 ;
        RECT 107.870 124.270 126.650 124.300 ;
        RECT 111.250 124.260 126.650 124.270 ;
        RECT 119.400 123.660 123.550 123.760 ;
        RECT 119.400 123.260 123.600 123.660 ;
        RECT 135.150 123.360 138.400 123.860 ;
        RECT 123.950 122.260 124.400 122.310 ;
        RECT 122.600 122.060 124.400 122.260 ;
        RECT 122.600 121.960 123.000 122.060 ;
        RECT 123.950 121.910 124.400 122.060 ;
        RECT 121.500 119.760 124.400 120.060 ;
        RECT 109.570 118.760 112.430 118.770 ;
        RECT 109.570 117.070 120.350 118.760 ;
        RECT 111.200 117.060 120.350 117.070 ;
        RECT 137.750 116.960 141.350 117.460 ;
        RECT 131.950 113.960 136.750 114.560 ;
        RECT 123.800 112.460 139.100 112.860 ;
        RECT 124.300 111.910 127.950 112.260 ;
        RECT 124.300 111.860 124.800 111.910 ;
        RECT 122.550 111.360 122.950 111.460 ;
        RECT 121.750 111.060 128.200 111.360 ;
        RECT 122.900 110.460 124.900 110.760 ;
        RECT 128.300 110.560 132.600 110.860 ;
        RECT 128.350 110.460 132.600 110.560 ;
        RECT 137.800 110.260 138.500 110.860 ;
        RECT 119.400 109.660 123.350 110.160 ;
        RECT 125.250 109.960 146.950 110.060 ;
        RECT 125.250 109.460 147.000 109.960 ;
        RECT 147.800 109.260 148.800 110.160 ;
        RECT 131.750 76.860 132.850 77.960 ;
      LAYER via2 ;
        RECT 49.100 194.500 50.500 196.200 ;
        RECT 145.950 176.760 146.750 179.260 ;
        RECT 90.300 174.000 91.300 174.900 ;
        RECT 96.500 171.100 97.300 171.900 ;
        RECT 153.750 160.460 155.150 162.060 ;
        RECT 147.050 151.960 148.850 152.960 ;
        RECT 129.260 149.620 130.660 151.720 ;
        RECT 128.360 142.820 129.660 145.020 ;
        RECT 103.300 130.500 104.100 131.300 ;
        RECT 103.300 127.500 104.100 128.300 ;
        RECT 88.100 125.800 88.900 126.600 ;
        RECT 1.000 124.300 2.400 125.400 ;
        RECT 137.850 110.260 138.450 110.860 ;
        RECT 119.550 109.660 120.050 110.160 ;
        RECT 147.850 109.260 148.750 110.160 ;
        RECT 131.850 76.960 132.750 77.860 ;
      LAYER met3 ;
        RECT 49.050 194.475 50.550 196.225 ;
        RECT 88.000 125.700 89.000 223.300 ;
        RECT 0.950 124.275 2.450 125.425 ;
        RECT 90.250 4.050 91.350 175.000 ;
        RECT 96.400 4.000 97.400 172.000 ;
        RECT 103.200 130.400 104.200 222.600 ;
        RECT 145.750 179.310 146.750 179.360 ;
        RECT 145.750 176.710 146.775 179.310 ;
        RECT 111.460 151.720 126.860 169.920 ;
        RECT 145.750 160.660 146.750 176.710 ;
        RECT 155.000 162.110 157.200 162.400 ;
        RECT 145.850 160.510 146.750 160.660 ;
        RECT 147.850 153.160 149.050 161.860 ;
        RECT 153.725 160.410 157.200 162.110 ;
        RECT 147.050 153.010 149.050 153.160 ;
        RECT 147.025 151.910 149.050 153.010 ;
        RECT 129.235 151.720 130.685 151.770 ;
        RECT 147.050 151.760 149.050 151.910 ;
        RECT 111.460 149.620 130.760 151.720 ;
        RECT 111.460 138.060 126.860 149.620 ;
        RECT 129.235 149.570 130.685 149.620 ;
        RECT 128.260 142.720 129.760 145.120 ;
        RECT 103.200 16.800 104.200 128.400 ;
        RECT 119.350 108.160 120.150 110.360 ;
        RECT 137.750 110.160 138.550 110.960 ;
        RECT 147.850 110.210 149.050 151.760 ;
        RECT 147.825 109.210 149.050 110.210 ;
        RECT 147.850 109.160 149.050 109.210 ;
        RECT 119.350 80.560 148.610 108.160 ;
        RECT 119.350 76.260 120.150 80.560 ;
        RECT 131.750 76.860 132.850 77.960 ;
        RECT 119.350 73.860 148.610 76.260 ;
        RECT 119.550 48.660 148.610 73.860 ;
        RECT 134.300 4.600 135.300 17.800 ;
        RECT 155.000 7.600 157.200 160.410 ;
      LAYER via3 ;
        RECT 88.100 222.400 88.900 223.100 ;
        RECT 49.100 194.500 50.500 196.200 ;
        RECT 103.300 221.700 104.100 222.500 ;
        RECT 1.000 124.300 2.400 125.400 ;
        RECT 90.300 4.200 91.300 5.100 ;
        RECT 145.850 160.560 146.750 162.160 ;
        RECT 147.950 160.460 148.950 161.760 ;
        RECT 153.750 160.460 155.150 162.060 ;
        RECT 128.360 142.820 129.660 145.020 ;
        RECT 111.600 138.160 126.720 138.480 ;
        RECT 137.850 110.260 138.450 110.860 ;
        RECT 119.650 80.700 119.970 108.020 ;
        RECT 131.850 76.960 132.750 77.860 ;
        RECT 119.650 48.800 119.970 76.120 ;
        RECT 103.300 16.900 104.100 17.700 ;
        RECT 134.400 16.900 135.200 17.700 ;
        RECT 96.500 4.100 97.300 4.900 ;
        RECT 155.200 7.800 157.000 9.600 ;
        RECT 134.400 4.700 135.200 5.500 ;
      LAYER met4 ;
        RECT 88.630 224.100 88.930 224.760 ;
        RECT 88.000 222.300 89.000 224.100 ;
        RECT 154.870 222.600 155.170 224.760 ;
        RECT 103.200 221.600 155.500 222.600 ;
        RECT 50.500 194.495 50.505 196.205 ;
        RECT 111.855 145.020 126.465 169.525 ;
        RECT 150.745 162.260 151.355 162.265 ;
        RECT 145.100 160.360 155.550 162.260 ;
        RECT 128.260 145.020 129.760 145.120 ;
        RECT 111.855 142.820 129.760 145.020 ;
        RECT 111.855 139.915 126.465 142.820 ;
        RECT 128.260 142.720 129.760 142.820 ;
        RECT 111.520 138.080 126.800 138.560 ;
        RECT 0.995 124.295 1.000 125.405 ;
        RECT 119.570 80.620 120.050 108.100 ;
        RECT 136.350 107.765 138.550 112.060 ;
        RECT 121.405 80.955 148.215 107.765 ;
        RECT 131.750 77.160 132.850 77.960 ;
        RECT 119.570 48.720 120.050 76.200 ;
        RECT 131.150 75.865 133.350 77.160 ;
        RECT 121.405 49.055 148.215 75.865 ;
        RECT 103.200 16.800 135.300 17.800 ;
        RECT 90.250 2.650 91.350 5.150 ;
        RECT 96.400 4.000 113.100 5.000 ;
        RECT 90.320 1.000 90.920 2.650 ;
        RECT 112.400 1.000 113.000 4.000 ;
        RECT 134.300 2.500 135.300 5.600 ;
        RECT 155.000 3.600 157.200 9.800 ;
        RECT 134.480 1.000 135.080 2.500 ;
        RECT 156.560 1.000 157.160 3.600 ;
  END
END tt_um_hugodg_temp_sensor
END LIBRARY

