MACRO device_without_rf
  CLASS BLOCK ;
  FOREIGN device_without_rf ;
  ORIGIN 0.310 12.900 ;
  SIZE 148.410 BY 50.600 ;
  PIN vd
    ANTENNAGATEAREA 8.000000 ;
    ANTENNADIFFAREA 49.667625 ;
    PORT
      LAYER met1 ;
        RECT 34.900 36.700 35.900 37.700 ;
    END
  END vd
  PIN gnd
    ANTENNAGATEAREA 18.000000 ;
    ANTENNADIFFAREA 39.573498 ;
    PORT
      LAYER met1 ;
        RECT -0.310 -9.780 0.690 -8.780 ;
    END
  END gnd
  PIN clk
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met1 ;
        RECT 65.390 -12.880 66.390 -11.880 ;
    END
  END clk
  PIN vpwr
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 1.764300 ;
    PORT
      LAYER met1 ;
        RECT 71.390 -12.880 72.390 -11.880 ;
    END
  END vpwr
  PIN ib
    ANTENNAGATEAREA 3.000000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met1 ;
        RECT 24.790 -12.880 25.790 -11.880 ;
    END
  END ib
  PIN out_buff
    ANTENNAGATEAREA 30.224998 ;
    ANTENNADIFFAREA 18.850000 ;
    PORT
      LAYER met1 ;
        RECT 68.290 -12.880 69.290 -11.880 ;
    END
  END out_buff
  PIN vts
    ANTENNAGATEAREA 4.225000 ;
    ANTENNADIFFAREA 12.156000 ;
    PORT
      LAYER met1 ;
        RECT 21.800 -12.900 22.800 -11.900 ;
    END
  END vts
  PIN out
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met1 ;
        RECT 70.090 -12.880 71.090 -11.880 ;
    END
  END out
  OBS
      LAYER nwell ;
        RECT 1.035 18.135 21.165 26.465 ;
        RECT 28.040 24.010 59.940 27.710 ;
        RECT 0.835 11.535 16.965 16.865 ;
      LAYER pwell ;
        RECT 0.000 0.800 16.960 10.400 ;
      LAYER nwell ;
        RECT 28.175 10.245 35.005 24.010 ;
      LAYER pwell ;
        RECT 36.540 20.010 52.500 23.910 ;
        RECT 36.540 17.810 43.440 20.010 ;
        RECT 43.540 17.810 52.500 20.010 ;
        RECT 36.540 12.910 52.500 17.810 ;
      LAYER nwell ;
        RECT 53.140 10.210 59.940 24.010 ;
      LAYER pwell ;
        RECT 71.800 10.600 87.760 29.700 ;
      LAYER nwell ;
        RECT 71.600 6.950 73.700 7.000 ;
        RECT 71.600 5.800 83.760 6.950 ;
        RECT 72.800 5.345 83.760 5.800 ;
      LAYER pwell ;
        RECT 77.505 4.825 78.435 5.045 ;
        RECT 81.155 4.825 83.510 5.055 ;
        RECT 72.995 4.145 83.510 4.825 ;
      LAYER nwell ;
        RECT 85.070 4.670 87.180 9.860 ;
      LAYER pwell ;
        RECT 73.135 3.955 73.305 4.145 ;
        RECT 85.070 1.320 87.180 4.420 ;
      LAYER li1 ;
        RECT 71.980 29.350 87.580 29.520 ;
        RECT 41.440 27.495 46.640 27.510 ;
        RECT 59.240 27.495 59.740 27.510 ;
        RECT 28.355 27.325 59.740 27.495 ;
        RECT 4.200 26.285 5.000 26.300 ;
        RECT 9.800 26.285 10.600 26.300 ;
        RECT 13.700 26.285 14.500 26.300 ;
        RECT 18.300 26.285 19.100 26.300 ;
        RECT 1.215 26.115 20.985 26.285 ;
        RECT 1.215 18.485 1.385 26.115 ;
        RECT 4.200 26.100 5.000 26.115 ;
        RECT 9.800 26.100 10.600 26.115 ;
        RECT 13.700 26.100 14.500 26.115 ;
        RECT 18.300 26.100 19.100 26.115 ;
        RECT 9.070 25.135 10.070 25.305 ;
        RECT 10.970 25.135 11.970 25.305 ;
        RECT 12.870 25.135 17.870 25.305 ;
        RECT 18.770 25.135 19.770 25.305 ;
        RECT 8.840 22.880 9.010 24.920 ;
        RECT 10.130 22.880 10.300 24.920 ;
        RECT 10.740 22.880 10.910 24.920 ;
        RECT 12.030 22.880 12.200 24.920 ;
        RECT 12.640 22.880 12.810 24.920 ;
        RECT 17.930 22.880 18.100 24.920 ;
        RECT 18.540 22.880 18.710 24.920 ;
        RECT 19.830 22.880 20.000 24.920 ;
        RECT 9.070 22.495 10.070 22.665 ;
        RECT 10.970 22.495 11.970 22.665 ;
        RECT 12.870 22.495 17.870 22.665 ;
        RECT 18.770 22.495 19.770 22.665 ;
        RECT 2.170 21.735 3.170 21.905 ;
        RECT 4.070 21.735 5.070 21.905 ;
        RECT 5.360 21.735 6.360 21.905 ;
        RECT 7.270 21.735 8.270 21.905 ;
        RECT 8.560 21.735 9.560 21.905 ;
        RECT 9.850 21.735 10.850 21.905 ;
        RECT 11.140 21.735 12.140 21.905 ;
        RECT 13.070 21.735 14.070 21.905 ;
        RECT 14.360 21.735 15.360 21.905 ;
        RECT 15.650 21.735 16.650 21.905 ;
        RECT 16.940 21.735 17.940 21.905 ;
        RECT 18.870 21.735 19.870 21.905 ;
        RECT 1.940 19.480 2.110 21.520 ;
        RECT 3.230 19.480 3.400 21.520 ;
        RECT 3.840 19.480 4.010 21.520 ;
        RECT 5.130 19.480 5.300 21.520 ;
        RECT 6.420 19.480 6.590 21.520 ;
        RECT 7.040 19.480 7.210 21.520 ;
        RECT 8.330 19.480 8.500 21.520 ;
        RECT 9.620 19.480 9.790 21.520 ;
        RECT 10.910 19.480 11.080 21.520 ;
        RECT 12.200 19.480 12.370 21.520 ;
        RECT 12.840 19.480 13.010 21.520 ;
        RECT 14.130 19.480 14.300 21.520 ;
        RECT 15.420 19.480 15.590 21.520 ;
        RECT 16.710 19.480 16.880 21.520 ;
        RECT 18.000 19.480 18.170 21.520 ;
        RECT 18.640 19.480 18.810 21.520 ;
        RECT 19.930 19.480 20.100 21.520 ;
        RECT 2.170 19.095 3.170 19.265 ;
        RECT 4.070 19.095 5.070 19.265 ;
        RECT 5.360 19.095 6.360 19.265 ;
        RECT 7.270 19.095 8.270 19.265 ;
        RECT 8.560 19.095 9.560 19.265 ;
        RECT 9.850 19.095 10.850 19.265 ;
        RECT 11.140 19.095 12.140 19.265 ;
        RECT 13.070 19.095 14.070 19.265 ;
        RECT 14.360 19.095 15.360 19.265 ;
        RECT 15.650 19.095 16.650 19.265 ;
        RECT 16.940 19.095 17.940 19.265 ;
        RECT 18.870 19.095 19.870 19.265 ;
        RECT 20.815 18.485 20.985 26.115 ;
        RECT 1.215 18.315 20.985 18.485 ;
        RECT 28.355 24.395 28.525 27.325 ;
        RECT 35.355 27.310 35.525 27.325 ;
        RECT 41.440 27.310 46.640 27.325 ;
        RECT 52.855 27.310 53.025 27.325 ;
        RECT 59.240 27.310 59.740 27.325 ;
        RECT 29.110 26.645 30.110 26.815 ;
        RECT 30.400 26.645 31.400 26.815 ;
        RECT 31.690 26.645 32.690 26.815 ;
        RECT 32.980 26.645 33.980 26.815 ;
        RECT 34.910 26.645 35.910 26.815 ;
        RECT 36.200 26.645 37.200 26.815 ;
        RECT 37.490 26.645 38.490 26.815 ;
        RECT 38.780 26.645 39.780 26.815 ;
        RECT 40.070 26.645 41.070 26.815 ;
        RECT 41.360 26.645 42.360 26.815 ;
        RECT 42.650 26.645 43.650 26.815 ;
        RECT 44.510 26.645 45.510 26.815 ;
        RECT 45.800 26.645 46.800 26.815 ;
        RECT 47.090 26.645 48.090 26.815 ;
        RECT 48.380 26.645 49.380 26.815 ;
        RECT 49.670 26.645 50.670 26.815 ;
        RECT 50.960 26.645 51.960 26.815 ;
        RECT 52.250 26.645 53.250 26.815 ;
        RECT 54.110 26.645 55.110 26.815 ;
        RECT 55.400 26.645 56.400 26.815 ;
        RECT 56.690 26.645 57.690 26.815 ;
        RECT 57.980 26.645 58.980 26.815 ;
        RECT 28.355 24.225 28.540 24.395 ;
        RECT 1.015 16.515 16.785 16.685 ;
        RECT 1.015 11.885 1.185 16.515 ;
        RECT 2.070 15.535 3.070 15.705 ;
        RECT 3.970 15.535 4.970 15.705 ;
        RECT 5.260 15.535 6.260 15.705 ;
        RECT 6.550 15.535 7.550 15.705 ;
        RECT 7.840 15.535 8.840 15.705 ;
        RECT 9.130 15.535 10.130 15.705 ;
        RECT 10.420 15.535 11.420 15.705 ;
        RECT 11.710 15.535 12.710 15.705 ;
        RECT 13.000 15.535 14.000 15.705 ;
        RECT 14.870 15.535 15.870 15.705 ;
        RECT 1.840 13.280 2.010 15.320 ;
        RECT 3.130 13.280 3.300 15.320 ;
        RECT 3.740 13.280 3.910 15.320 ;
        RECT 5.030 13.280 5.200 15.320 ;
        RECT 6.320 13.280 6.490 15.320 ;
        RECT 7.610 13.280 7.780 15.320 ;
        RECT 8.900 13.280 9.070 15.320 ;
        RECT 10.190 13.280 10.360 15.320 ;
        RECT 11.480 13.280 11.650 15.320 ;
        RECT 12.770 13.280 12.940 15.320 ;
        RECT 14.060 13.280 14.230 15.320 ;
        RECT 14.640 13.280 14.810 15.320 ;
        RECT 15.930 13.280 16.100 15.320 ;
        RECT 16.615 15.200 16.785 16.515 ;
        RECT 16.400 14.700 16.800 15.200 ;
        RECT 2.070 12.895 3.070 13.065 ;
        RECT 3.970 12.895 4.970 13.065 ;
        RECT 5.260 12.895 6.260 13.065 ;
        RECT 6.550 12.895 7.550 13.065 ;
        RECT 7.840 12.895 8.840 13.065 ;
        RECT 9.130 12.895 10.130 13.065 ;
        RECT 10.420 12.895 11.420 13.065 ;
        RECT 11.710 12.895 12.710 13.065 ;
        RECT 13.000 12.895 14.000 13.065 ;
        RECT 14.870 12.895 15.870 13.065 ;
        RECT 16.615 11.885 16.785 14.700 ;
        RECT 1.015 11.715 16.785 11.885 ;
        RECT 28.355 10.595 28.525 24.225 ;
        RECT 28.880 11.390 29.050 26.430 ;
        RECT 30.170 11.390 30.340 26.430 ;
        RECT 31.460 11.390 31.630 26.430 ;
        RECT 32.750 11.390 32.920 26.430 ;
        RECT 34.040 11.390 34.210 26.430 ;
        RECT 34.680 25.390 34.850 26.430 ;
        RECT 35.970 25.390 36.140 26.430 ;
        RECT 37.260 25.390 37.430 26.430 ;
        RECT 38.550 25.390 38.720 26.430 ;
        RECT 39.840 25.390 40.010 26.430 ;
        RECT 41.130 25.390 41.300 26.430 ;
        RECT 42.420 25.390 42.590 26.430 ;
        RECT 43.710 25.390 43.880 26.430 ;
        RECT 44.280 25.390 44.450 26.430 ;
        RECT 45.570 25.390 45.740 26.430 ;
        RECT 46.860 25.390 47.030 26.430 ;
        RECT 48.150 25.390 48.320 26.430 ;
        RECT 49.440 25.390 49.610 26.430 ;
        RECT 50.730 25.390 50.900 26.430 ;
        RECT 52.020 25.390 52.190 26.430 ;
        RECT 53.310 25.390 53.480 26.430 ;
        RECT 34.910 25.005 35.910 25.175 ;
        RECT 36.200 25.005 37.200 25.175 ;
        RECT 37.490 25.005 38.490 25.175 ;
        RECT 38.780 25.005 39.780 25.175 ;
        RECT 40.070 25.005 41.070 25.175 ;
        RECT 41.360 25.005 42.360 25.175 ;
        RECT 42.650 25.005 43.650 25.175 ;
        RECT 44.510 25.005 45.530 25.175 ;
        RECT 45.800 25.005 46.820 25.175 ;
        RECT 47.090 25.005 48.110 25.175 ;
        RECT 48.380 25.005 49.400 25.175 ;
        RECT 49.670 25.005 50.690 25.175 ;
        RECT 50.960 25.005 51.960 25.175 ;
        RECT 52.250 25.005 53.270 25.175 ;
        RECT 34.740 24.395 36.040 24.410 ;
        RECT 53.355 24.395 53.525 24.410 ;
        RECT 34.640 24.225 53.525 24.395 ;
        RECT 34.640 24.210 36.040 24.225 ;
        RECT 34.640 23.825 34.825 24.210 ;
        RECT 29.110 11.005 30.110 11.175 ;
        RECT 30.400 11.005 31.400 11.175 ;
        RECT 31.690 11.005 32.690 11.175 ;
        RECT 32.980 11.005 33.980 11.175 ;
        RECT 34.655 10.595 34.825 23.825 ;
        RECT 36.720 23.660 52.320 23.830 ;
        RECT 36.720 13.260 36.890 23.660 ;
        RECT 43.840 23.240 44.170 23.410 ;
        RECT 44.800 23.240 45.130 23.410 ;
        RECT 43.200 21.530 43.370 23.070 ;
        RECT 43.680 21.530 43.850 23.070 ;
        RECT 44.160 21.530 44.330 23.070 ;
        RECT 44.640 21.530 44.810 23.070 ;
        RECT 45.120 21.530 45.290 23.070 ;
        RECT 43.360 21.190 43.690 21.360 ;
        RECT 44.320 21.190 44.650 21.360 ;
        RECT 38.330 19.640 39.330 19.810 ;
        RECT 39.620 19.640 40.620 19.810 ;
        RECT 40.910 19.640 41.910 19.810 ;
        RECT 42.200 19.640 43.200 19.810 ;
        RECT 38.100 18.430 38.270 19.470 ;
        RECT 39.390 18.430 39.560 19.470 ;
        RECT 40.680 18.430 40.850 19.470 ;
        RECT 41.970 18.430 42.140 19.470 ;
        RECT 43.260 18.430 43.430 19.470 ;
        RECT 44.130 19.340 45.130 19.510 ;
        RECT 45.420 19.340 46.420 19.510 ;
        RECT 46.710 19.340 47.710 19.510 ;
        RECT 48.000 19.340 49.000 19.510 ;
        RECT 49.290 19.340 50.290 19.510 ;
        RECT 50.580 19.340 51.580 19.510 ;
        RECT 38.330 18.090 39.330 18.260 ;
        RECT 39.620 18.090 40.620 18.260 ;
        RECT 40.910 18.090 41.910 18.260 ;
        RECT 42.200 18.090 43.200 18.260 ;
        RECT 43.900 14.130 44.070 19.170 ;
        RECT 45.190 14.130 45.360 19.170 ;
        RECT 46.480 14.130 46.650 19.170 ;
        RECT 47.770 14.130 47.940 19.170 ;
        RECT 49.060 14.130 49.230 19.170 ;
        RECT 50.350 14.130 50.520 19.170 ;
        RECT 51.640 14.130 51.810 19.170 ;
        RECT 44.130 13.790 45.130 13.960 ;
        RECT 45.420 13.790 46.420 13.960 ;
        RECT 46.710 13.790 47.710 13.960 ;
        RECT 48.000 13.790 49.000 13.960 ;
        RECT 49.290 13.790 50.290 13.960 ;
        RECT 50.580 13.790 51.580 13.960 ;
        RECT 40.540 13.260 41.040 13.410 ;
        RECT 47.640 13.260 48.140 13.410 ;
        RECT 52.150 13.260 52.320 23.660 ;
        RECT 36.720 13.090 52.320 13.260 ;
        RECT 40.540 13.010 41.040 13.090 ;
        RECT 47.640 13.010 48.140 13.090 ;
        RECT 28.355 10.425 34.825 10.595 ;
        RECT 53.355 10.595 53.525 24.225 ;
        RECT 53.880 11.390 54.050 26.430 ;
        RECT 55.170 11.390 55.340 26.430 ;
        RECT 56.460 11.390 56.630 26.430 ;
        RECT 57.750 11.390 57.920 26.430 ;
        RECT 59.040 11.390 59.210 26.430 ;
        RECT 59.555 24.395 59.725 27.310 ;
        RECT 59.540 24.225 59.725 24.395 ;
        RECT 54.110 11.005 55.110 11.175 ;
        RECT 55.400 11.005 56.400 11.175 ;
        RECT 56.690 11.005 57.690 11.175 ;
        RECT 57.980 11.005 58.980 11.175 ;
        RECT 59.555 10.595 59.725 24.225 ;
        RECT 71.980 10.950 72.150 29.350 ;
        RECT 72.750 26.600 73.100 28.760 ;
        RECT 73.580 26.600 73.930 28.760 ;
        RECT 74.410 26.600 74.760 28.760 ;
        RECT 75.240 26.600 75.590 28.760 ;
        RECT 76.070 26.600 76.420 28.760 ;
        RECT 76.900 26.600 77.250 28.760 ;
        RECT 77.730 26.600 78.080 28.760 ;
        RECT 78.560 26.600 78.910 28.760 ;
        RECT 80.120 26.600 80.470 28.760 ;
        RECT 80.950 26.600 81.300 28.760 ;
        RECT 81.780 26.600 82.130 28.760 ;
        RECT 82.610 26.600 82.960 28.760 ;
        RECT 83.440 26.600 83.790 28.760 ;
        RECT 84.270 26.600 84.620 28.760 ;
        RECT 85.100 26.600 85.450 28.760 ;
        RECT 85.930 26.600 86.280 28.760 ;
        RECT 72.750 19.940 73.100 22.100 ;
        RECT 73.580 19.940 73.930 22.100 ;
        RECT 74.410 19.940 74.760 22.100 ;
        RECT 75.240 19.940 75.590 22.100 ;
        RECT 76.070 19.940 76.420 22.100 ;
        RECT 76.900 19.940 77.250 22.100 ;
        RECT 77.730 19.940 78.080 22.100 ;
        RECT 78.560 19.940 78.910 22.100 ;
        RECT 80.120 19.940 80.470 22.100 ;
        RECT 80.950 19.940 81.300 22.100 ;
        RECT 81.780 19.940 82.130 22.100 ;
        RECT 82.610 19.940 82.960 22.100 ;
        RECT 83.440 19.940 83.790 22.100 ;
        RECT 84.270 19.940 84.620 22.100 ;
        RECT 85.100 19.940 85.450 22.100 ;
        RECT 85.930 19.940 86.280 22.100 ;
        RECT 73.000 15.760 73.350 17.920 ;
        RECT 73.830 15.760 74.180 17.920 ;
        RECT 74.660 15.760 75.010 17.920 ;
        RECT 75.490 15.760 75.840 17.920 ;
        RECT 76.320 15.760 76.670 17.920 ;
        RECT 77.150 15.760 77.500 17.920 ;
        RECT 77.980 15.760 78.330 17.920 ;
        RECT 78.810 15.760 79.160 17.920 ;
        RECT 73.000 11.600 73.350 13.760 ;
        RECT 73.830 11.600 74.180 13.760 ;
        RECT 74.660 11.600 75.010 13.760 ;
        RECT 75.490 11.600 75.840 13.760 ;
        RECT 76.320 11.600 76.670 13.760 ;
        RECT 77.150 11.600 77.500 13.760 ;
        RECT 77.980 11.600 78.330 13.760 ;
        RECT 78.810 11.600 79.160 13.760 ;
        RECT 80.100 10.950 80.700 11.000 ;
        RECT 87.410 10.950 87.580 29.350 ;
        RECT 71.980 10.780 87.580 10.950 ;
        RECT 53.355 10.425 59.725 10.595 ;
        RECT 0.180 10.050 16.780 10.220 ;
        RECT 0.180 1.150 0.350 10.050 ;
        RECT 1.090 9.550 2.090 9.720 ;
        RECT 2.990 9.550 3.990 9.720 ;
        RECT 4.890 9.550 5.890 9.720 ;
        RECT 6.790 9.550 7.790 9.720 ;
        RECT 8.690 9.550 9.690 9.720 ;
        RECT 10.590 9.550 11.590 9.720 ;
        RECT 12.490 9.550 13.490 9.720 ;
        RECT 14.390 9.550 15.390 9.720 ;
        RECT 0.860 8.340 1.030 9.380 ;
        RECT 2.150 8.340 2.320 9.380 ;
        RECT 2.760 8.340 2.930 9.380 ;
        RECT 4.050 8.340 4.220 9.380 ;
        RECT 4.660 8.340 4.830 9.380 ;
        RECT 5.950 8.340 6.120 9.380 ;
        RECT 6.560 8.340 6.730 9.380 ;
        RECT 7.850 8.340 8.020 9.380 ;
        RECT 8.460 8.340 8.630 9.380 ;
        RECT 9.750 8.340 9.920 9.380 ;
        RECT 10.360 8.340 10.530 9.380 ;
        RECT 11.650 8.340 11.820 9.380 ;
        RECT 12.260 8.340 12.430 9.380 ;
        RECT 13.550 8.340 13.720 9.380 ;
        RECT 14.160 8.340 14.330 9.380 ;
        RECT 15.450 8.340 15.620 9.380 ;
        RECT 1.090 8.000 2.090 8.170 ;
        RECT 2.990 8.000 3.990 8.170 ;
        RECT 4.890 8.000 5.890 8.170 ;
        RECT 6.790 8.000 7.790 8.170 ;
        RECT 8.690 8.000 9.690 8.170 ;
        RECT 10.590 8.000 11.590 8.170 ;
        RECT 12.490 8.000 13.490 8.170 ;
        RECT 14.390 8.000 15.390 8.170 ;
        RECT 1.090 7.460 2.090 7.630 ;
        RECT 2.990 7.460 3.990 7.630 ;
        RECT 4.890 7.460 5.890 7.630 ;
        RECT 6.790 7.460 7.790 7.630 ;
        RECT 8.690 7.460 9.690 7.630 ;
        RECT 10.590 7.460 11.590 7.630 ;
        RECT 12.490 7.460 13.490 7.630 ;
        RECT 14.390 7.460 15.390 7.630 ;
        RECT 0.860 6.250 1.030 7.290 ;
        RECT 2.150 6.250 2.320 7.290 ;
        RECT 2.760 6.250 2.930 7.290 ;
        RECT 4.050 6.250 4.220 7.290 ;
        RECT 4.660 6.250 4.830 7.290 ;
        RECT 5.950 6.250 6.120 7.290 ;
        RECT 6.560 6.250 6.730 7.290 ;
        RECT 7.850 6.250 8.020 7.290 ;
        RECT 8.460 6.250 8.630 7.290 ;
        RECT 9.750 6.250 9.920 7.290 ;
        RECT 10.360 6.250 10.530 7.290 ;
        RECT 11.650 6.250 11.820 7.290 ;
        RECT 12.260 6.250 12.430 7.290 ;
        RECT 13.550 6.250 13.720 7.290 ;
        RECT 14.160 6.250 14.330 7.290 ;
        RECT 15.450 6.250 15.620 7.290 ;
        RECT 1.090 5.910 2.090 6.080 ;
        RECT 2.990 5.910 3.990 6.080 ;
        RECT 4.890 5.910 5.890 6.080 ;
        RECT 6.790 5.910 7.790 6.080 ;
        RECT 8.690 5.910 9.690 6.080 ;
        RECT 10.590 5.910 11.590 6.080 ;
        RECT 12.490 5.910 13.490 6.080 ;
        RECT 14.390 5.910 15.390 6.080 ;
        RECT 1.090 5.370 2.090 5.540 ;
        RECT 2.990 5.370 3.990 5.540 ;
        RECT 4.890 5.370 5.890 5.540 ;
        RECT 6.790 5.370 7.790 5.540 ;
        RECT 8.690 5.370 9.690 5.540 ;
        RECT 10.590 5.370 11.590 5.540 ;
        RECT 12.490 5.370 13.490 5.540 ;
        RECT 14.390 5.370 15.390 5.540 ;
        RECT 0.860 4.160 1.030 5.200 ;
        RECT 2.150 4.160 2.320 5.200 ;
        RECT 2.760 4.160 2.930 5.200 ;
        RECT 4.050 4.160 4.220 5.200 ;
        RECT 4.660 4.160 4.830 5.200 ;
        RECT 5.950 4.160 6.120 5.200 ;
        RECT 6.560 4.160 6.730 5.200 ;
        RECT 7.850 4.160 8.020 5.200 ;
        RECT 8.460 4.160 8.630 5.200 ;
        RECT 9.750 4.160 9.920 5.200 ;
        RECT 10.360 4.160 10.530 5.200 ;
        RECT 11.650 4.160 11.820 5.200 ;
        RECT 12.260 4.160 12.430 5.200 ;
        RECT 13.550 4.160 13.720 5.200 ;
        RECT 14.160 4.160 14.330 5.200 ;
        RECT 15.450 4.160 15.620 5.200 ;
        RECT 1.090 3.820 2.090 3.990 ;
        RECT 2.990 3.820 3.990 3.990 ;
        RECT 4.890 3.820 5.890 3.990 ;
        RECT 6.790 3.820 7.790 3.990 ;
        RECT 8.690 3.820 9.690 3.990 ;
        RECT 10.590 3.820 11.590 3.990 ;
        RECT 12.490 3.820 13.490 3.990 ;
        RECT 14.390 3.820 15.390 3.990 ;
        RECT 1.090 3.280 2.090 3.450 ;
        RECT 2.990 3.280 3.990 3.450 ;
        RECT 4.890 3.280 5.890 3.450 ;
        RECT 6.790 3.280 7.790 3.450 ;
        RECT 8.690 3.280 9.690 3.450 ;
        RECT 10.590 3.280 11.590 3.450 ;
        RECT 12.490 3.280 13.490 3.450 ;
        RECT 14.390 3.280 15.390 3.450 ;
        RECT 0.860 2.070 1.030 3.110 ;
        RECT 2.150 2.070 2.320 3.110 ;
        RECT 2.760 2.070 2.930 3.110 ;
        RECT 4.050 2.070 4.220 3.110 ;
        RECT 4.660 2.070 4.830 3.110 ;
        RECT 5.950 2.070 6.120 3.110 ;
        RECT 6.560 2.070 6.730 3.110 ;
        RECT 7.850 2.070 8.020 3.110 ;
        RECT 8.460 2.070 8.630 3.110 ;
        RECT 9.750 2.070 9.920 3.110 ;
        RECT 10.360 2.070 10.530 3.110 ;
        RECT 11.650 2.070 11.820 3.110 ;
        RECT 12.260 2.070 12.430 3.110 ;
        RECT 13.550 2.070 13.720 3.110 ;
        RECT 14.160 2.070 14.330 3.110 ;
        RECT 15.450 2.070 15.620 3.110 ;
        RECT 1.090 1.730 2.090 1.900 ;
        RECT 2.990 1.730 3.990 1.900 ;
        RECT 4.890 1.730 5.890 1.900 ;
        RECT 6.790 1.730 7.790 1.900 ;
        RECT 8.690 1.730 9.690 1.900 ;
        RECT 10.590 1.730 11.590 1.900 ;
        RECT 12.490 1.730 13.490 1.900 ;
        RECT 14.390 1.730 15.390 1.900 ;
        RECT 1.100 1.150 2.200 1.200 ;
        RECT 5.500 1.150 6.600 1.200 ;
        RECT 10.100 1.150 11.200 1.200 ;
        RECT 14.300 1.150 15.400 1.200 ;
        RECT 16.610 1.150 16.780 10.050 ;
        RECT 85.250 9.510 87.000 9.680 ;
        RECT 72.990 6.675 83.570 6.845 ;
        RECT 72.100 6.100 72.600 6.550 ;
        RECT 73.080 6.005 73.335 6.505 ;
        RECT 73.505 6.175 73.835 6.675 ;
        RECT 73.080 5.835 73.830 6.005 ;
        RECT 73.080 5.015 73.430 5.665 ;
        RECT 73.600 4.845 73.830 5.835 ;
        RECT 73.080 4.675 73.830 4.845 ;
        RECT 73.080 4.385 73.335 4.675 ;
        RECT 73.505 4.125 73.835 4.505 ;
        RECT 74.005 4.385 74.175 6.505 ;
        RECT 74.345 5.705 74.670 6.490 ;
        RECT 74.840 6.215 75.090 6.675 ;
        RECT 75.260 6.175 75.510 6.505 ;
        RECT 75.725 6.175 76.405 6.505 ;
        RECT 75.260 6.045 75.430 6.175 ;
        RECT 75.035 5.875 75.430 6.045 ;
        RECT 74.405 4.655 74.865 5.705 ;
        RECT 75.035 4.515 75.205 5.875 ;
        RECT 75.600 5.615 76.065 6.005 ;
        RECT 75.375 4.805 75.725 5.425 ;
        RECT 75.895 5.025 76.065 5.615 ;
        RECT 76.235 5.395 76.405 6.175 ;
        RECT 76.575 6.075 76.745 6.415 ;
        RECT 76.980 6.245 77.310 6.675 ;
        RECT 77.480 6.075 77.650 6.415 ;
        RECT 77.945 6.215 78.315 6.675 ;
        RECT 76.575 5.905 77.650 6.075 ;
        RECT 78.485 6.045 78.655 6.505 ;
        RECT 78.890 6.165 79.760 6.505 ;
        RECT 79.930 6.215 80.180 6.675 ;
        RECT 78.095 5.875 78.655 6.045 ;
        RECT 78.095 5.735 78.265 5.875 ;
        RECT 76.765 5.565 78.265 5.735 ;
        RECT 78.960 5.705 79.420 5.995 ;
        RECT 76.235 5.225 77.925 5.395 ;
        RECT 75.895 4.805 76.250 5.025 ;
        RECT 76.420 4.515 76.590 5.225 ;
        RECT 76.795 4.805 77.585 5.055 ;
        RECT 77.755 5.045 77.925 5.225 ;
        RECT 78.095 4.875 78.265 5.565 ;
        RECT 74.535 4.125 74.865 4.485 ;
        RECT 75.035 4.345 75.530 4.515 ;
        RECT 75.735 4.345 76.590 4.515 ;
        RECT 77.465 4.125 77.795 4.585 ;
        RECT 78.005 4.485 78.265 4.875 ;
        RECT 78.455 5.695 79.420 5.705 ;
        RECT 79.590 5.785 79.760 6.165 ;
        RECT 80.350 6.125 80.520 6.415 ;
        RECT 80.700 6.295 81.420 6.675 ;
        RECT 80.350 5.955 81.150 6.125 ;
        RECT 78.455 5.535 79.130 5.695 ;
        RECT 79.590 5.615 80.810 5.785 ;
        RECT 78.455 4.745 78.665 5.535 ;
        RECT 79.590 5.525 79.760 5.615 ;
        RECT 78.835 4.745 79.185 5.365 ;
        RECT 79.355 5.355 79.760 5.525 ;
        RECT 79.355 4.575 79.525 5.355 ;
        RECT 79.695 4.905 79.915 5.185 ;
        RECT 80.095 5.075 80.635 5.445 ;
        RECT 80.980 5.365 81.150 5.955 ;
        RECT 81.590 5.495 81.995 6.505 ;
        RECT 80.980 5.335 81.425 5.365 ;
        RECT 79.695 4.735 80.225 4.905 ;
        RECT 78.005 4.315 78.355 4.485 ;
        RECT 78.575 4.295 79.525 4.575 ;
        RECT 79.695 4.125 79.885 4.565 ;
        RECT 80.055 4.505 80.225 4.735 ;
        RECT 80.395 4.675 80.635 5.075 ;
        RECT 80.805 5.035 81.425 5.335 ;
        RECT 80.805 4.860 81.130 5.035 ;
        RECT 80.805 4.505 81.125 4.860 ;
        RECT 80.055 4.335 81.125 4.505 ;
        RECT 81.325 4.125 81.495 4.810 ;
        RECT 81.665 4.800 81.995 5.495 ;
        RECT 82.185 5.365 82.515 6.465 ;
        RECT 82.750 5.535 82.920 6.675 ;
        RECT 83.170 5.485 83.425 6.365 ;
        RECT 82.185 5.035 83.045 5.365 ;
        RECT 83.215 5.300 83.425 5.485 ;
        RECT 83.215 5.100 83.450 5.300 ;
        RECT 81.665 4.500 82.000 4.800 ;
        RECT 81.665 4.315 81.995 4.500 ;
        RECT 82.185 4.385 82.435 5.035 ;
        RECT 83.215 4.835 83.425 5.100 ;
        RECT 85.250 5.020 85.420 9.510 ;
        RECT 85.960 9.000 86.290 9.170 ;
        RECT 85.820 5.745 85.990 8.785 ;
        RECT 86.260 5.745 86.430 8.785 ;
        RECT 86.830 8.700 87.000 9.510 ;
        RECT 86.800 5.900 87.000 8.700 ;
        RECT 85.960 5.360 86.290 5.530 ;
        RECT 86.830 5.020 87.000 5.900 ;
        RECT 85.250 4.850 87.000 5.020 ;
        RECT 82.750 4.125 82.920 4.720 ;
        RECT 83.170 4.305 83.425 4.835 ;
        RECT 72.990 3.955 83.570 4.125 ;
        RECT 85.250 4.070 87.000 4.240 ;
        RECT 85.250 1.670 85.420 4.070 ;
        RECT 85.960 3.560 86.290 3.730 ;
        RECT 85.820 2.350 85.990 3.390 ;
        RECT 86.260 2.350 86.430 3.390 ;
        RECT 86.830 3.200 87.000 4.070 ;
        RECT 86.800 2.400 87.000 3.200 ;
        RECT 85.960 2.010 86.290 2.180 ;
        RECT 86.830 1.670 87.000 2.400 ;
        RECT 85.250 1.500 87.000 1.670 ;
        RECT 0.180 0.980 16.780 1.150 ;
      LAYER mcon ;
        RECT 9.150 25.135 9.990 25.305 ;
        RECT 11.050 25.135 11.890 25.305 ;
        RECT 12.950 25.135 17.790 25.305 ;
        RECT 18.850 25.135 19.690 25.305 ;
        RECT 8.840 23.815 9.010 24.755 ;
        RECT 10.130 23.815 10.300 24.755 ;
        RECT 10.740 22.960 10.910 24.840 ;
        RECT 12.030 22.960 12.200 24.840 ;
        RECT 12.640 22.960 12.810 24.840 ;
        RECT 17.930 22.960 18.100 24.840 ;
        RECT 18.540 23.815 18.710 24.755 ;
        RECT 19.830 23.815 20.000 24.755 ;
        RECT 9.150 22.495 9.990 22.665 ;
        RECT 11.050 22.495 11.890 22.665 ;
        RECT 12.950 22.495 17.790 22.665 ;
        RECT 18.850 22.495 19.690 22.665 ;
        RECT 2.250 21.735 3.090 21.905 ;
        RECT 4.150 21.735 4.990 21.905 ;
        RECT 5.440 21.735 6.280 21.905 ;
        RECT 7.350 21.735 8.190 21.905 ;
        RECT 8.640 21.735 9.480 21.905 ;
        RECT 9.930 21.735 10.770 21.905 ;
        RECT 11.220 21.735 12.060 21.905 ;
        RECT 13.150 21.735 13.990 21.905 ;
        RECT 14.440 21.735 15.280 21.905 ;
        RECT 15.730 21.735 16.570 21.905 ;
        RECT 17.020 21.735 17.860 21.905 ;
        RECT 18.950 21.735 19.790 21.905 ;
        RECT 1.940 20.415 2.110 21.355 ;
        RECT 3.230 20.415 3.400 21.355 ;
        RECT 3.840 19.645 4.010 20.585 ;
        RECT 5.130 20.415 5.300 21.355 ;
        RECT 6.420 19.645 6.590 20.585 ;
        RECT 7.040 19.645 7.210 20.585 ;
        RECT 8.330 20.415 8.500 21.355 ;
        RECT 9.620 19.645 9.790 20.585 ;
        RECT 10.910 20.415 11.080 21.355 ;
        RECT 12.200 19.645 12.370 20.585 ;
        RECT 12.840 19.645 13.010 20.585 ;
        RECT 14.130 20.415 14.300 21.355 ;
        RECT 15.420 19.645 15.590 20.585 ;
        RECT 16.710 20.415 16.880 21.355 ;
        RECT 18.000 19.645 18.170 20.585 ;
        RECT 18.640 19.645 18.810 20.585 ;
        RECT 19.930 19.645 20.100 20.585 ;
        RECT 2.250 19.095 3.090 19.265 ;
        RECT 4.150 19.095 4.990 19.265 ;
        RECT 5.440 19.095 6.280 19.265 ;
        RECT 7.350 19.095 8.190 19.265 ;
        RECT 8.640 19.095 9.480 19.265 ;
        RECT 9.930 19.095 10.770 19.265 ;
        RECT 11.220 19.095 12.060 19.265 ;
        RECT 13.150 19.095 13.990 19.265 ;
        RECT 14.440 19.095 15.280 19.265 ;
        RECT 15.730 19.095 16.570 19.265 ;
        RECT 17.020 19.095 17.860 19.265 ;
        RECT 18.950 19.095 19.790 19.265 ;
        RECT 30.480 26.645 31.320 26.815 ;
        RECT 31.770 26.645 32.610 26.815 ;
        RECT 36.280 26.645 37.120 26.815 ;
        RECT 51.040 26.645 51.880 26.815 ;
        RECT 55.480 26.645 56.320 26.815 ;
        RECT 56.770 26.645 57.610 26.815 ;
        RECT 2.150 15.535 2.990 15.705 ;
        RECT 4.050 15.535 4.890 15.705 ;
        RECT 5.340 15.535 6.180 15.705 ;
        RECT 6.630 15.535 7.470 15.705 ;
        RECT 7.920 15.535 8.760 15.705 ;
        RECT 9.210 15.535 10.050 15.705 ;
        RECT 10.500 15.535 11.340 15.705 ;
        RECT 11.790 15.535 12.630 15.705 ;
        RECT 13.080 15.535 13.920 15.705 ;
        RECT 14.950 15.535 15.790 15.705 ;
        RECT 1.840 14.215 2.010 15.155 ;
        RECT 3.130 14.215 3.300 15.155 ;
        RECT 3.740 13.445 3.910 14.385 ;
        RECT 5.030 14.215 5.200 15.155 ;
        RECT 6.320 13.445 6.490 14.385 ;
        RECT 7.610 14.215 7.780 15.155 ;
        RECT 8.900 13.445 9.070 14.385 ;
        RECT 10.190 14.215 10.360 15.155 ;
        RECT 11.480 13.445 11.650 14.385 ;
        RECT 12.770 14.215 12.940 15.155 ;
        RECT 14.060 13.445 14.230 14.385 ;
        RECT 14.640 14.215 14.810 15.155 ;
        RECT 15.930 14.215 16.100 15.155 ;
        RECT 16.400 14.700 16.800 15.200 ;
        RECT 2.150 12.895 2.990 13.065 ;
        RECT 4.050 12.895 4.890 13.065 ;
        RECT 5.340 12.895 6.180 13.065 ;
        RECT 6.630 12.895 7.470 13.065 ;
        RECT 7.920 12.895 8.760 13.065 ;
        RECT 9.210 12.895 10.050 13.065 ;
        RECT 10.500 12.895 11.340 13.065 ;
        RECT 11.790 12.895 12.630 13.065 ;
        RECT 13.080 12.895 13.920 13.065 ;
        RECT 14.950 12.895 15.790 13.065 ;
        RECT 28.880 18.825 29.050 26.265 ;
        RECT 30.170 11.555 30.340 18.995 ;
        RECT 31.460 18.825 31.630 26.265 ;
        RECT 32.750 11.555 32.920 18.995 ;
        RECT 34.040 18.825 34.210 26.265 ;
        RECT 34.680 25.555 34.850 25.995 ;
        RECT 35.970 25.825 36.140 26.265 ;
        RECT 37.260 25.555 37.430 25.995 ;
        RECT 38.550 25.825 38.720 26.265 ;
        RECT 39.840 25.555 40.010 25.995 ;
        RECT 41.130 25.825 41.300 26.265 ;
        RECT 42.420 25.555 42.590 25.995 ;
        RECT 43.710 25.825 43.880 26.265 ;
        RECT 44.280 25.555 44.450 25.995 ;
        RECT 45.570 25.825 45.740 26.265 ;
        RECT 46.860 25.555 47.030 25.995 ;
        RECT 48.150 25.825 48.320 26.265 ;
        RECT 49.440 25.555 49.610 25.995 ;
        RECT 50.730 25.825 50.900 26.265 ;
        RECT 52.020 25.555 52.190 25.995 ;
        RECT 53.310 25.825 53.480 26.265 ;
        RECT 34.990 25.005 35.830 25.175 ;
        RECT 36.280 25.005 37.120 25.175 ;
        RECT 37.570 25.005 38.410 25.175 ;
        RECT 38.860 25.005 39.700 25.175 ;
        RECT 40.150 25.005 40.990 25.175 ;
        RECT 41.440 25.005 42.280 25.175 ;
        RECT 42.730 25.005 43.570 25.175 ;
        RECT 44.690 25.005 45.530 25.175 ;
        RECT 45.980 25.005 46.820 25.175 ;
        RECT 47.270 25.005 48.110 25.175 ;
        RECT 48.560 25.005 49.400 25.175 ;
        RECT 49.850 25.005 50.690 25.175 ;
        RECT 51.040 25.005 51.880 25.175 ;
        RECT 52.330 25.005 53.270 25.175 ;
        RECT 29.190 11.005 30.030 11.175 ;
        RECT 33.060 11.005 33.900 11.175 ;
        RECT 43.920 23.240 44.090 23.410 ;
        RECT 44.880 23.240 45.050 23.410 ;
        RECT 43.200 21.695 43.370 22.385 ;
        RECT 43.680 22.215 43.850 22.905 ;
        RECT 44.160 21.695 44.330 22.385 ;
        RECT 44.640 22.215 44.810 22.905 ;
        RECT 45.120 21.695 45.290 22.385 ;
        RECT 43.440 21.190 43.610 21.360 ;
        RECT 44.400 21.190 44.570 21.360 ;
        RECT 38.410 19.640 39.250 19.810 ;
        RECT 39.700 19.640 40.540 19.810 ;
        RECT 40.990 19.640 41.830 19.810 ;
        RECT 42.280 19.640 43.120 19.810 ;
        RECT 38.100 18.595 38.270 19.035 ;
        RECT 39.390 18.865 39.560 19.305 ;
        RECT 40.680 18.595 40.850 19.035 ;
        RECT 41.970 18.865 42.140 19.305 ;
        RECT 44.210 19.340 45.050 19.510 ;
        RECT 45.500 19.340 46.340 19.510 ;
        RECT 46.790 19.340 47.630 19.510 ;
        RECT 48.080 19.340 48.920 19.510 ;
        RECT 49.370 19.340 50.210 19.510 ;
        RECT 50.660 19.340 51.500 19.510 ;
        RECT 43.260 18.595 43.430 19.035 ;
        RECT 38.410 18.090 39.250 18.260 ;
        RECT 39.700 18.090 40.540 18.260 ;
        RECT 40.990 18.090 41.830 18.260 ;
        RECT 42.280 18.090 43.120 18.260 ;
        RECT 43.900 16.565 44.070 19.005 ;
        RECT 45.190 14.295 45.360 16.735 ;
        RECT 46.480 16.565 46.650 19.005 ;
        RECT 47.770 14.295 47.940 16.735 ;
        RECT 49.060 16.565 49.230 19.005 ;
        RECT 50.350 14.295 50.520 16.735 ;
        RECT 51.640 16.565 51.810 19.005 ;
        RECT 44.210 13.790 45.050 13.960 ;
        RECT 45.500 13.790 46.340 13.960 ;
        RECT 46.790 13.790 47.630 13.960 ;
        RECT 48.080 13.790 48.920 13.960 ;
        RECT 49.370 13.790 50.210 13.960 ;
        RECT 50.660 13.790 51.500 13.960 ;
        RECT 53.880 18.825 54.050 26.265 ;
        RECT 55.170 11.555 55.340 18.995 ;
        RECT 56.460 18.825 56.630 26.265 ;
        RECT 57.750 11.555 57.920 18.995 ;
        RECT 59.040 18.825 59.210 26.265 ;
        RECT 54.190 11.005 55.030 11.175 ;
        RECT 58.060 11.005 58.900 11.175 ;
        RECT 72.830 26.685 73.020 28.670 ;
        RECT 73.660 26.685 73.850 28.670 ;
        RECT 74.490 26.685 74.680 28.670 ;
        RECT 75.320 26.685 75.510 28.670 ;
        RECT 76.150 26.685 76.340 28.670 ;
        RECT 76.980 26.685 77.170 28.670 ;
        RECT 77.810 26.685 78.000 28.670 ;
        RECT 78.640 26.685 78.830 28.670 ;
        RECT 80.200 26.685 80.390 28.670 ;
        RECT 81.030 26.685 81.220 28.670 ;
        RECT 81.860 26.685 82.050 28.670 ;
        RECT 82.690 26.685 82.880 28.670 ;
        RECT 83.520 26.685 83.710 28.670 ;
        RECT 84.350 26.685 84.540 28.670 ;
        RECT 85.180 26.685 85.370 28.670 ;
        RECT 86.010 26.685 86.200 28.670 ;
        RECT 72.830 20.030 73.020 22.015 ;
        RECT 73.660 20.030 73.850 22.015 ;
        RECT 74.490 20.030 74.680 22.015 ;
        RECT 75.320 20.030 75.510 22.015 ;
        RECT 76.150 20.030 76.340 22.015 ;
        RECT 76.980 20.030 77.170 22.015 ;
        RECT 77.810 20.030 78.000 22.015 ;
        RECT 78.640 20.030 78.830 22.015 ;
        RECT 80.200 20.030 80.390 22.015 ;
        RECT 81.030 20.030 81.220 22.015 ;
        RECT 81.860 20.030 82.050 22.015 ;
        RECT 82.690 20.030 82.880 22.015 ;
        RECT 83.520 20.030 83.710 22.015 ;
        RECT 84.350 20.030 84.540 22.015 ;
        RECT 85.180 20.030 85.370 22.015 ;
        RECT 86.010 20.030 86.200 22.015 ;
        RECT 73.080 15.845 73.270 17.830 ;
        RECT 73.910 15.845 74.100 17.830 ;
        RECT 74.740 15.845 74.930 17.830 ;
        RECT 75.570 15.845 75.760 17.830 ;
        RECT 76.400 15.845 76.590 17.830 ;
        RECT 77.230 15.845 77.420 17.830 ;
        RECT 78.060 15.845 78.250 17.830 ;
        RECT 78.890 15.845 79.080 17.830 ;
        RECT 73.080 11.690 73.270 13.675 ;
        RECT 73.910 11.690 74.100 13.675 ;
        RECT 74.740 11.690 74.930 13.675 ;
        RECT 75.570 11.690 75.760 13.675 ;
        RECT 76.400 11.690 76.590 13.675 ;
        RECT 77.230 11.690 77.420 13.675 ;
        RECT 78.060 11.690 78.250 13.675 ;
        RECT 78.890 11.690 79.080 13.675 ;
        RECT 1.170 9.550 2.010 9.720 ;
        RECT 3.070 9.550 3.910 9.720 ;
        RECT 4.970 9.550 5.810 9.720 ;
        RECT 6.870 9.550 7.710 9.720 ;
        RECT 8.770 9.550 9.610 9.720 ;
        RECT 10.670 9.550 11.510 9.720 ;
        RECT 12.570 9.550 13.410 9.720 ;
        RECT 14.470 9.550 15.310 9.720 ;
        RECT 0.860 8.420 1.030 9.300 ;
        RECT 2.150 8.420 2.320 9.300 ;
        RECT 2.760 8.420 2.930 9.300 ;
        RECT 4.050 8.420 4.220 9.300 ;
        RECT 4.660 8.420 4.830 9.300 ;
        RECT 5.950 8.420 6.120 9.300 ;
        RECT 6.560 8.420 6.730 9.300 ;
        RECT 7.850 8.420 8.020 9.300 ;
        RECT 8.460 8.420 8.630 9.300 ;
        RECT 9.750 8.420 9.920 9.300 ;
        RECT 10.360 8.420 10.530 9.300 ;
        RECT 11.650 8.420 11.820 9.300 ;
        RECT 12.260 8.420 12.430 9.300 ;
        RECT 13.550 8.420 13.720 9.300 ;
        RECT 14.160 8.420 14.330 9.300 ;
        RECT 15.450 8.420 15.620 9.300 ;
        RECT 1.170 8.000 2.010 8.170 ;
        RECT 3.070 8.000 3.910 8.170 ;
        RECT 4.970 8.000 5.810 8.170 ;
        RECT 6.870 8.000 7.710 8.170 ;
        RECT 8.770 8.000 9.610 8.170 ;
        RECT 10.670 8.000 11.510 8.170 ;
        RECT 12.570 8.000 13.410 8.170 ;
        RECT 14.470 8.000 15.310 8.170 ;
        RECT 1.170 7.460 2.010 7.630 ;
        RECT 3.070 7.460 3.910 7.630 ;
        RECT 4.970 7.460 5.810 7.630 ;
        RECT 6.870 7.460 7.710 7.630 ;
        RECT 8.770 7.460 9.610 7.630 ;
        RECT 10.670 7.460 11.510 7.630 ;
        RECT 12.570 7.460 13.410 7.630 ;
        RECT 14.470 7.460 15.310 7.630 ;
        RECT 0.860 6.330 1.030 7.210 ;
        RECT 2.150 6.330 2.320 7.210 ;
        RECT 2.760 6.330 2.930 7.210 ;
        RECT 4.050 6.330 4.220 7.210 ;
        RECT 4.660 6.330 4.830 7.210 ;
        RECT 5.950 6.330 6.120 7.210 ;
        RECT 6.560 6.330 6.730 7.210 ;
        RECT 7.850 6.330 8.020 7.210 ;
        RECT 8.460 6.330 8.630 7.210 ;
        RECT 9.750 6.330 9.920 7.210 ;
        RECT 10.360 6.330 10.530 7.210 ;
        RECT 11.650 6.330 11.820 7.210 ;
        RECT 12.260 6.330 12.430 7.210 ;
        RECT 13.550 6.330 13.720 7.210 ;
        RECT 14.160 6.330 14.330 7.210 ;
        RECT 15.450 6.330 15.620 7.210 ;
        RECT 1.170 5.910 2.010 6.080 ;
        RECT 3.070 5.910 3.910 6.080 ;
        RECT 4.970 5.910 5.810 6.080 ;
        RECT 6.870 5.910 7.710 6.080 ;
        RECT 8.770 5.910 9.610 6.080 ;
        RECT 10.670 5.910 11.510 6.080 ;
        RECT 12.570 5.910 13.410 6.080 ;
        RECT 14.470 5.910 15.310 6.080 ;
        RECT 1.170 5.370 2.010 5.540 ;
        RECT 3.070 5.370 3.910 5.540 ;
        RECT 4.970 5.370 5.810 5.540 ;
        RECT 6.870 5.370 7.710 5.540 ;
        RECT 8.770 5.370 9.610 5.540 ;
        RECT 10.670 5.370 11.510 5.540 ;
        RECT 12.570 5.370 13.410 5.540 ;
        RECT 14.470 5.370 15.310 5.540 ;
        RECT 0.860 4.240 1.030 5.120 ;
        RECT 2.150 4.240 2.320 5.120 ;
        RECT 2.760 4.240 2.930 5.120 ;
        RECT 4.050 4.240 4.220 5.120 ;
        RECT 4.660 4.240 4.830 5.120 ;
        RECT 5.950 4.240 6.120 5.120 ;
        RECT 6.560 4.240 6.730 5.120 ;
        RECT 7.850 4.240 8.020 5.120 ;
        RECT 8.460 4.240 8.630 5.120 ;
        RECT 9.750 4.240 9.920 5.120 ;
        RECT 10.360 4.240 10.530 5.120 ;
        RECT 11.650 4.240 11.820 5.120 ;
        RECT 12.260 4.240 12.430 5.120 ;
        RECT 13.550 4.240 13.720 5.120 ;
        RECT 14.160 4.240 14.330 5.120 ;
        RECT 15.450 4.240 15.620 5.120 ;
        RECT 1.170 3.820 2.010 3.990 ;
        RECT 3.070 3.820 3.910 3.990 ;
        RECT 4.970 3.820 5.810 3.990 ;
        RECT 6.870 3.820 7.710 3.990 ;
        RECT 8.770 3.820 9.610 3.990 ;
        RECT 10.670 3.820 11.510 3.990 ;
        RECT 12.570 3.820 13.410 3.990 ;
        RECT 14.470 3.820 15.310 3.990 ;
        RECT 1.170 3.280 2.010 3.450 ;
        RECT 3.070 3.280 3.910 3.450 ;
        RECT 4.970 3.280 5.810 3.450 ;
        RECT 6.870 3.280 7.710 3.450 ;
        RECT 8.770 3.280 9.610 3.450 ;
        RECT 10.670 3.280 11.510 3.450 ;
        RECT 12.570 3.280 13.410 3.450 ;
        RECT 14.470 3.280 15.310 3.450 ;
        RECT 0.860 2.150 1.030 3.030 ;
        RECT 2.150 2.150 2.320 3.030 ;
        RECT 2.760 2.150 2.930 3.030 ;
        RECT 4.050 2.150 4.220 3.030 ;
        RECT 4.660 2.150 4.830 3.030 ;
        RECT 5.950 2.150 6.120 3.030 ;
        RECT 6.560 2.150 6.730 3.030 ;
        RECT 7.850 2.150 8.020 3.030 ;
        RECT 8.460 2.150 8.630 3.030 ;
        RECT 9.750 2.150 9.920 3.030 ;
        RECT 10.360 2.150 10.530 3.030 ;
        RECT 11.650 2.150 11.820 3.030 ;
        RECT 12.260 2.150 12.430 3.030 ;
        RECT 13.550 2.150 13.720 3.030 ;
        RECT 14.160 2.150 14.330 3.030 ;
        RECT 15.450 2.150 15.620 3.030 ;
        RECT 1.170 1.730 2.010 1.900 ;
        RECT 3.070 1.730 3.910 1.900 ;
        RECT 4.970 1.730 5.810 1.900 ;
        RECT 6.870 1.730 7.710 1.900 ;
        RECT 8.770 1.730 9.610 1.900 ;
        RECT 10.670 1.730 11.510 1.900 ;
        RECT 12.570 1.730 13.410 1.900 ;
        RECT 14.470 1.730 15.310 1.900 ;
        RECT 1.100 1.000 2.200 1.200 ;
        RECT 5.500 1.000 6.600 1.200 ;
        RECT 10.100 1.000 11.200 1.200 ;
        RECT 14.300 1.000 15.400 1.200 ;
        RECT 73.135 6.675 73.305 6.845 ;
        RECT 73.595 6.675 73.765 6.845 ;
        RECT 74.055 6.675 74.225 6.845 ;
        RECT 74.515 6.675 74.685 6.845 ;
        RECT 74.975 6.675 75.145 6.845 ;
        RECT 75.435 6.675 75.605 6.845 ;
        RECT 75.895 6.675 76.065 6.845 ;
        RECT 76.355 6.675 76.525 6.845 ;
        RECT 76.815 6.675 76.985 6.845 ;
        RECT 77.275 6.675 77.445 6.845 ;
        RECT 77.735 6.675 77.905 6.845 ;
        RECT 78.195 6.675 78.365 6.845 ;
        RECT 78.655 6.675 78.825 6.845 ;
        RECT 79.115 6.675 79.285 6.845 ;
        RECT 79.575 6.675 79.745 6.845 ;
        RECT 80.035 6.675 80.205 6.845 ;
        RECT 80.495 6.675 80.665 6.845 ;
        RECT 80.955 6.675 81.125 6.845 ;
        RECT 81.415 6.675 81.585 6.845 ;
        RECT 81.875 6.675 82.045 6.845 ;
        RECT 82.335 6.675 82.505 6.845 ;
        RECT 82.795 6.675 82.965 6.845 ;
        RECT 83.255 6.675 83.425 6.845 ;
        RECT 72.150 6.250 72.500 6.500 ;
        RECT 73.100 5.100 73.300 5.400 ;
        RECT 73.600 5.145 73.770 5.315 ;
        RECT 74.005 5.825 74.175 5.995 ;
        RECT 74.500 4.750 74.800 4.950 ;
        RECT 75.895 5.825 76.065 5.995 ;
        RECT 75.435 5.145 75.605 5.315 ;
        RECT 79.015 5.825 79.185 5.995 ;
        RECT 77.155 4.805 77.325 4.975 ;
        RECT 79.015 5.145 79.185 5.315 ;
        RECT 80.095 5.120 80.265 5.290 ;
        RECT 80.395 4.805 80.565 4.975 ;
        RECT 83.250 5.100 83.450 5.300 ;
        RECT 81.700 4.500 82.000 4.800 ;
        RECT 86.040 9.000 86.210 9.170 ;
        RECT 85.820 5.825 85.990 8.705 ;
        RECT 86.260 5.825 86.430 8.705 ;
        RECT 86.800 5.900 87.000 8.700 ;
        RECT 86.040 5.360 86.210 5.530 ;
        RECT 73.135 3.955 73.305 4.125 ;
        RECT 73.595 3.955 73.765 4.125 ;
        RECT 74.055 3.955 74.225 4.125 ;
        RECT 74.515 3.955 74.685 4.125 ;
        RECT 74.975 3.955 75.145 4.125 ;
        RECT 75.435 3.955 75.605 4.125 ;
        RECT 75.895 3.955 76.065 4.125 ;
        RECT 76.355 3.955 76.525 4.125 ;
        RECT 76.815 3.955 76.985 4.125 ;
        RECT 77.275 3.955 77.445 4.125 ;
        RECT 77.735 3.955 77.905 4.125 ;
        RECT 78.195 3.955 78.365 4.125 ;
        RECT 78.655 3.955 78.825 4.125 ;
        RECT 79.115 3.955 79.285 4.125 ;
        RECT 79.575 3.955 79.745 4.125 ;
        RECT 80.035 3.955 80.205 4.125 ;
        RECT 80.495 3.955 80.665 4.125 ;
        RECT 80.955 3.955 81.125 4.125 ;
        RECT 81.415 3.955 81.585 4.125 ;
        RECT 81.875 3.955 82.045 4.125 ;
        RECT 82.335 3.955 82.505 4.125 ;
        RECT 82.795 3.955 82.965 4.125 ;
        RECT 83.255 3.955 83.425 4.125 ;
        RECT 86.040 3.560 86.210 3.730 ;
        RECT 85.820 2.430 85.990 3.310 ;
        RECT 86.260 2.430 86.430 3.310 ;
        RECT 86.800 2.400 87.000 3.200 ;
        RECT 86.040 2.010 86.210 2.180 ;
      LAYER met1 ;
        RECT 34.700 36.700 34.900 37.700 ;
        RECT 35.900 36.700 36.300 37.700 ;
        RECT 34.700 36.000 36.300 36.700 ;
        RECT 34.500 34.300 36.500 36.000 ;
        RECT 43.750 28.710 44.850 29.500 ;
        RECT 31.340 27.710 42.340 27.810 ;
        RECT 43.740 27.710 44.850 28.710 ;
        RECT 72.800 28.700 73.050 28.730 ;
        RECT 73.630 28.700 73.880 28.730 ;
        RECT 1.600 27.000 21.200 27.500 ;
        RECT 31.340 27.110 56.840 27.710 ;
        RECT 1.550 26.500 21.200 27.000 ;
        RECT 30.420 26.810 31.380 26.845 ;
        RECT 31.710 26.810 32.670 26.845 ;
        RECT 36.220 26.810 37.180 26.845 ;
        RECT 29.140 26.615 37.180 26.810 ;
        RECT 29.140 26.610 37.140 26.615 ;
        RECT 50.940 26.610 58.940 26.910 ;
        RECT 4.200 26.330 5.000 26.500 ;
        RECT 9.800 26.330 10.600 26.500 ;
        RECT 13.700 26.330 14.500 26.500 ;
        RECT 18.300 26.330 19.100 26.500 ;
        RECT 4.140 26.070 5.060 26.330 ;
        RECT 9.740 26.070 10.660 26.330 ;
        RECT 13.640 26.070 14.560 26.330 ;
        RECT 18.240 26.070 19.160 26.330 ;
        RECT 9.100 25.335 10.200 25.400 ;
        RECT 9.090 25.300 10.200 25.335 ;
        RECT 9.000 24.815 10.200 25.300 ;
        RECT 10.990 25.105 11.950 25.335 ;
        RECT 12.890 25.105 17.850 25.335 ;
        RECT 18.790 25.300 19.750 25.335 ;
        RECT 18.790 25.200 19.900 25.300 ;
        RECT 8.810 24.800 10.330 24.815 ;
        RECT 10.710 24.800 10.940 24.900 ;
        RECT 7.950 24.200 11.000 24.800 ;
        RECT 8.810 23.755 9.040 24.200 ;
        RECT 10.100 23.755 10.330 24.200 ;
        RECT 10.710 22.900 10.940 24.200 ;
        RECT 12.000 24.000 12.230 24.900 ;
        RECT 11.750 22.900 12.250 24.000 ;
        RECT 12.610 23.800 12.840 24.900 ;
        RECT 17.900 24.800 18.130 24.900 ;
        RECT 18.600 24.815 19.900 25.200 ;
        RECT 18.510 24.800 20.030 24.815 ;
        RECT 17.900 24.200 20.750 24.800 ;
        RECT 17.900 24.100 20.100 24.200 ;
        RECT 12.600 23.700 16.900 23.800 ;
        RECT 12.600 23.100 16.950 23.700 ;
        RECT 12.610 22.900 12.840 23.100 ;
        RECT 17.900 22.900 18.130 24.100 ;
        RECT 18.510 23.755 18.740 24.100 ;
        RECT 19.800 23.755 20.030 24.100 ;
        RECT 11.000 22.695 13.650 22.700 ;
        RECT 9.090 22.465 10.050 22.695 ;
        RECT 10.990 22.500 17.850 22.695 ;
        RECT 10.990 22.465 11.950 22.500 ;
        RECT 12.890 22.465 17.850 22.500 ;
        RECT 18.790 22.465 19.750 22.695 ;
        RECT 13.050 22.400 13.650 22.465 ;
        RECT 2.190 21.900 3.150 21.935 ;
        RECT 2.190 21.705 3.200 21.900 ;
        RECT 4.090 21.705 5.050 21.935 ;
        RECT 5.380 21.705 6.340 21.935 ;
        RECT 7.290 21.705 8.250 21.935 ;
        RECT 8.580 21.705 9.540 21.935 ;
        RECT 9.870 21.705 10.830 21.935 ;
        RECT 11.160 21.705 12.120 21.935 ;
        RECT 13.090 21.705 14.050 21.935 ;
        RECT 14.380 21.705 15.340 21.935 ;
        RECT 15.670 21.705 16.630 21.935 ;
        RECT 16.960 21.705 17.920 21.935 ;
        RECT 18.890 21.705 19.850 21.935 ;
        RECT 2.200 21.500 3.200 21.705 ;
        RECT 1.550 21.415 5.300 21.500 ;
        RECT 1.550 21.100 5.330 21.415 ;
        RECT 1.910 20.355 2.140 21.100 ;
        RECT 3.200 20.355 3.430 21.100 ;
        RECT 3.810 20.100 4.040 20.645 ;
        RECT 5.100 20.355 5.330 21.100 ;
        RECT 8.300 21.000 12.500 21.500 ;
        RECT 14.100 21.400 14.330 21.415 ;
        RECT 16.680 21.400 16.910 21.415 ;
        RECT 6.390 20.100 6.620 20.645 ;
        RECT 3.800 19.585 6.620 20.100 ;
        RECT 7.010 20.000 7.240 20.645 ;
        RECT 8.300 20.355 8.530 21.000 ;
        RECT 9.590 20.000 9.820 20.645 ;
        RECT 10.880 20.355 11.110 21.000 ;
        RECT 14.100 20.900 16.910 21.400 ;
        RECT 12.170 20.000 12.400 20.645 ;
        RECT 12.810 20.000 13.040 20.645 ;
        RECT 14.100 20.355 14.330 20.900 ;
        RECT 15.390 20.000 15.620 20.645 ;
        RECT 16.680 20.355 16.910 20.900 ;
        RECT 17.970 20.000 18.200 20.645 ;
        RECT 18.610 20.000 18.840 20.645 ;
        RECT 19.900 20.000 20.130 20.645 ;
        RECT 3.800 19.300 6.600 19.585 ;
        RECT 7.000 19.500 20.200 20.000 ;
        RECT 3.800 19.295 12.100 19.300 ;
        RECT 13.050 19.295 17.900 19.300 ;
        RECT 18.900 19.295 19.800 19.500 ;
        RECT 28.850 19.310 29.080 26.325 ;
        RECT 31.430 25.610 31.660 26.325 ;
        RECT 31.290 24.410 31.890 25.610 ;
        RECT 2.190 19.065 3.150 19.295 ;
        RECT 3.800 19.200 12.120 19.295 ;
        RECT 4.090 19.065 12.120 19.200 ;
        RECT 13.050 19.100 17.920 19.295 ;
        RECT 13.050 19.065 14.050 19.100 ;
        RECT 14.380 19.065 15.340 19.100 ;
        RECT 15.670 19.065 16.630 19.100 ;
        RECT 16.960 19.065 17.920 19.100 ;
        RECT 18.890 19.065 19.850 19.295 ;
        RECT 4.100 19.000 12.100 19.065 ;
        RECT 13.050 19.000 13.650 19.065 ;
        RECT 28.840 19.055 30.240 19.310 ;
        RECT 28.840 18.410 30.370 19.055 ;
        RECT 31.430 18.765 31.660 24.410 ;
        RECT 34.010 19.310 34.240 26.325 ;
        RECT 35.940 26.210 41.490 26.410 ;
        RECT 34.740 26.055 36.170 26.210 ;
        RECT 34.650 25.765 36.170 26.055 ;
        RECT 34.650 25.495 36.040 25.765 ;
        RECT 37.230 25.610 37.460 26.055 ;
        RECT 38.520 25.765 38.750 26.210 ;
        RECT 39.810 25.610 40.040 26.055 ;
        RECT 40.890 26.010 41.490 26.210 ;
        RECT 42.540 26.325 43.840 26.410 ;
        RECT 45.640 26.325 50.940 26.410 ;
        RECT 42.540 26.055 43.910 26.325 ;
        RECT 45.540 26.210 50.940 26.325 ;
        RECT 53.280 26.310 53.510 26.325 ;
        RECT 44.440 26.055 45.990 26.210 ;
        RECT 41.100 25.765 41.330 26.010 ;
        RECT 42.390 25.910 43.910 26.055 ;
        RECT 42.290 25.765 43.910 25.910 ;
        RECT 44.250 25.810 45.990 26.055 ;
        RECT 46.830 26.010 47.060 26.055 ;
        RECT 44.250 25.765 45.770 25.810 ;
        RECT 42.290 25.610 43.840 25.765 ;
        RECT 34.740 25.010 36.040 25.495 ;
        RECT 37.140 25.410 43.840 25.610 ;
        RECT 44.250 25.510 45.740 25.765 ;
        RECT 46.690 25.610 47.190 26.010 ;
        RECT 48.120 25.765 48.350 26.210 ;
        RECT 49.410 25.610 49.640 26.055 ;
        RECT 50.700 25.765 50.930 26.210 ;
        RECT 51.990 26.010 52.220 26.055 ;
        RECT 52.740 26.010 53.540 26.310 ;
        RECT 51.990 25.810 53.540 26.010 ;
        RECT 51.990 25.765 53.510 25.810 ;
        RECT 51.990 25.610 53.440 25.765 ;
        RECT 44.250 25.495 46.040 25.510 ;
        RECT 41.340 25.210 42.340 25.410 ;
        RECT 36.240 25.205 42.340 25.210 ;
        RECT 36.220 25.010 42.340 25.205 ;
        RECT 42.540 25.010 43.840 25.410 ;
        RECT 44.440 25.210 46.040 25.495 ;
        RECT 46.690 25.410 53.440 25.610 ;
        RECT 44.440 25.205 51.840 25.210 ;
        RECT 44.440 25.010 51.940 25.205 ;
        RECT 52.240 25.110 53.440 25.410 ;
        RECT 34.930 24.975 35.890 25.010 ;
        RECT 36.220 24.975 37.180 25.010 ;
        RECT 37.510 24.975 38.470 25.010 ;
        RECT 38.800 24.975 39.760 25.010 ;
        RECT 40.090 24.975 41.050 25.010 ;
        RECT 41.380 24.975 42.340 25.010 ;
        RECT 42.670 24.975 43.630 25.010 ;
        RECT 44.630 24.975 45.590 25.010 ;
        RECT 45.920 24.975 46.880 25.010 ;
        RECT 47.210 24.975 48.170 25.010 ;
        RECT 48.500 24.975 49.460 25.010 ;
        RECT 49.790 24.975 50.750 25.010 ;
        RECT 50.980 24.975 51.940 25.010 ;
        RECT 52.270 25.010 53.440 25.110 ;
        RECT 52.270 24.975 53.330 25.010 ;
        RECT 43.790 23.710 53.090 24.110 ;
        RECT 43.790 23.210 44.290 23.510 ;
        RECT 44.840 23.440 45.140 23.510 ;
        RECT 44.820 23.310 45.140 23.440 ;
        RECT 44.740 23.010 45.240 23.310 ;
        RECT 42.290 22.965 43.740 23.010 ;
        RECT 44.740 22.965 45.990 23.010 ;
        RECT 42.290 22.610 43.880 22.965 ;
        RECT 43.140 22.155 43.880 22.610 ;
        RECT 44.610 22.610 45.990 22.965 ;
        RECT 44.610 22.445 45.240 22.610 ;
        RECT 43.140 21.610 43.740 22.155 ;
        RECT 44.130 22.010 44.360 22.445 ;
        RECT 44.610 22.155 45.320 22.445 ;
        RECT 43.990 21.610 44.390 22.010 ;
        RECT 44.740 21.910 45.320 22.155 ;
        RECT 45.090 21.635 45.320 21.910 ;
        RECT 43.340 21.110 43.740 21.610 ;
        RECT 44.340 21.310 44.640 21.410 ;
        RECT 45.490 21.310 45.890 21.410 ;
        RECT 44.340 21.110 45.940 21.310 ;
        RECT 35.190 20.510 45.940 20.810 ;
        RECT 41.890 20.010 44.390 20.310 ;
        RECT 38.350 19.610 39.310 19.840 ;
        RECT 39.640 19.610 40.600 19.840 ;
        RECT 40.930 19.610 41.890 19.840 ;
        RECT 42.220 19.810 43.180 19.840 ;
        RECT 42.220 19.610 43.340 19.810 ;
        RECT 32.740 19.055 34.240 19.310 ;
        RECT 38.440 19.110 39.140 19.610 ;
        RECT 42.340 19.410 43.340 19.610 ;
        RECT 45.540 19.540 50.240 19.610 ;
        RECT 44.150 19.510 45.110 19.540 ;
        RECT 42.040 19.365 43.340 19.410 ;
        RECT 39.360 19.110 39.590 19.365 ;
        RECT 41.940 19.310 43.340 19.365 ;
        RECT 32.720 18.765 34.240 19.055 ;
        RECT 20.200 17.700 21.850 17.800 ;
        RECT 13.050 17.100 21.850 17.700 ;
        RECT 13.100 17.000 21.850 17.100 ;
        RECT 20.200 16.800 21.850 17.000 ;
        RECT 1.900 15.215 3.200 15.800 ;
        RECT 3.990 15.505 4.950 15.735 ;
        RECT 5.280 15.505 6.240 15.735 ;
        RECT 6.570 15.505 7.530 15.735 ;
        RECT 7.860 15.505 8.820 15.735 ;
        RECT 9.150 15.505 10.110 15.735 ;
        RECT 10.440 15.505 11.400 15.735 ;
        RECT 11.730 15.505 12.690 15.735 ;
        RECT 13.020 15.505 13.980 15.735 ;
        RECT 14.800 15.215 15.900 15.800 ;
        RECT 30.140 15.710 30.370 18.410 ;
        RECT 32.720 18.410 34.140 18.765 ;
        RECT 38.040 18.710 39.990 19.110 ;
        RECT 41.890 19.095 43.340 19.310 ;
        RECT 43.940 19.310 45.110 19.510 ;
        RECT 45.440 19.310 50.270 19.540 ;
        RECT 50.600 19.510 51.560 19.540 ;
        RECT 50.600 19.310 51.740 19.510 ;
        RECT 40.650 19.010 40.880 19.095 ;
        RECT 38.070 18.535 38.300 18.710 ;
        RECT 32.720 15.710 32.950 18.410 ;
        RECT 38.440 18.290 39.140 18.710 ;
        RECT 39.540 18.310 39.940 18.710 ;
        RECT 40.490 18.510 41.090 19.010 ;
        RECT 41.890 18.810 43.460 19.095 ;
        RECT 43.940 19.065 45.040 19.310 ;
        RECT 41.940 18.805 43.460 18.810 ;
        RECT 42.040 18.710 43.460 18.805 ;
        RECT 42.340 18.535 43.460 18.710 ;
        RECT 43.870 18.810 45.040 19.065 ;
        RECT 45.540 19.065 46.540 19.310 ;
        RECT 50.640 19.065 51.740 19.310 ;
        RECT 53.850 19.210 54.080 26.325 ;
        RECT 56.430 26.210 56.660 26.325 ;
        RECT 56.290 23.410 56.690 26.210 ;
        RECT 38.350 18.060 39.310 18.290 ;
        RECT 39.540 18.110 41.940 18.310 ;
        RECT 42.340 18.290 43.340 18.535 ;
        RECT 42.220 18.110 43.340 18.290 ;
        RECT 39.640 18.060 40.600 18.110 ;
        RECT 40.930 18.060 41.890 18.110 ;
        RECT 42.220 18.060 43.180 18.110 ;
        RECT 43.870 16.810 44.100 18.810 ;
        RECT 45.540 18.510 46.680 19.065 ;
        RECT 44.240 18.010 46.680 18.510 ;
        RECT 43.840 16.795 45.340 16.810 ;
        RECT 43.840 16.210 45.390 16.795 ;
        RECT 46.450 16.505 46.680 18.010 ;
        RECT 49.030 17.910 49.260 19.065 ;
        RECT 50.640 18.610 51.840 19.065 ;
        RECT 49.030 17.410 51.340 17.910 ;
        RECT 1.810 15.200 3.330 15.215 ;
        RECT 5.000 15.200 5.230 15.215 ;
        RECT 7.580 15.200 7.810 15.215 ;
        RECT 10.160 15.200 10.390 15.215 ;
        RECT 12.740 15.200 12.970 15.215 ;
        RECT 14.610 15.200 16.130 15.215 ;
        RECT 16.370 15.200 16.830 15.260 ;
        RECT 20.200 15.200 27.800 15.500 ;
        RECT 1.800 14.700 27.800 15.200 ;
        RECT 1.810 14.155 2.040 14.700 ;
        RECT 3.100 14.155 3.330 14.700 ;
        RECT 3.710 14.000 3.940 14.445 ;
        RECT 5.000 14.155 5.230 14.700 ;
        RECT 6.290 14.000 6.520 14.445 ;
        RECT 7.580 14.155 7.810 14.700 ;
        RECT 8.870 14.000 9.100 14.445 ;
        RECT 10.160 14.155 10.390 14.700 ;
        RECT 11.450 14.000 11.680 14.445 ;
        RECT 12.740 14.155 12.970 14.700 ;
        RECT 14.030 14.000 14.260 14.445 ;
        RECT 14.610 14.155 14.840 14.700 ;
        RECT 15.900 14.155 16.130 14.700 ;
        RECT 16.370 14.640 16.830 14.700 ;
        RECT 20.200 14.500 27.800 14.700 ;
        RECT 30.140 15.210 44.690 15.710 ;
        RECT 45.160 15.610 45.390 16.210 ;
        RECT 47.740 15.610 47.970 16.795 ;
        RECT 49.030 16.505 49.260 17.410 ;
        RECT 51.610 16.810 51.840 18.610 ;
        RECT 53.840 19.055 55.340 19.210 ;
        RECT 53.840 18.310 55.370 19.055 ;
        RECT 56.430 18.765 56.660 23.410 ;
        RECT 59.010 19.210 59.240 26.325 ;
        RECT 60.100 26.100 72.400 27.100 ;
        RECT 72.700 26.700 73.880 28.700 ;
        RECT 72.800 26.625 73.050 26.700 ;
        RECT 73.630 26.625 73.880 26.700 ;
        RECT 74.460 28.700 74.710 28.730 ;
        RECT 75.290 28.700 75.540 28.730 ;
        RECT 76.120 28.700 76.370 28.730 ;
        RECT 76.950 28.700 77.200 28.730 ;
        RECT 74.460 26.700 75.600 28.700 ;
        RECT 76.100 26.700 77.200 28.700 ;
        RECT 74.460 26.625 74.710 26.700 ;
        RECT 75.290 26.625 75.540 26.700 ;
        RECT 76.120 26.625 76.370 26.700 ;
        RECT 76.950 26.625 77.200 26.700 ;
        RECT 77.780 28.700 78.030 28.730 ;
        RECT 78.610 28.700 78.860 28.730 ;
        RECT 80.170 28.700 80.420 28.730 ;
        RECT 81.000 28.700 81.250 28.730 ;
        RECT 81.830 28.700 82.080 28.730 ;
        RECT 82.660 28.700 82.910 28.730 ;
        RECT 83.490 28.700 83.740 28.730 ;
        RECT 84.320 28.700 84.570 28.730 ;
        RECT 85.150 28.700 85.400 28.730 ;
        RECT 85.980 28.700 86.230 28.730 ;
        RECT 77.780 26.700 78.900 28.700 ;
        RECT 80.170 26.700 81.300 28.700 ;
        RECT 81.830 26.700 83.000 28.700 ;
        RECT 83.490 26.700 84.600 28.700 ;
        RECT 85.150 26.700 86.300 28.700 ;
        RECT 86.550 28.500 87.700 29.400 ;
        RECT 86.700 28.400 87.700 28.500 ;
        RECT 86.700 27.600 87.300 28.400 ;
        RECT 86.700 27.200 87.350 27.600 ;
        RECT 77.780 26.625 78.030 26.700 ;
        RECT 78.610 26.625 78.860 26.700 ;
        RECT 80.170 26.625 80.420 26.700 ;
        RECT 81.000 26.625 81.250 26.700 ;
        RECT 81.830 26.625 82.080 26.700 ;
        RECT 82.660 26.625 82.910 26.700 ;
        RECT 83.490 26.625 83.740 26.700 ;
        RECT 84.320 26.625 84.570 26.700 ;
        RECT 85.150 26.625 85.400 26.700 ;
        RECT 85.980 26.625 86.230 26.700 ;
        RECT 72.500 21.700 73.100 22.100 ;
        RECT 73.630 22.000 73.880 22.075 ;
        RECT 74.460 22.000 74.710 22.075 ;
        RECT 71.500 20.700 73.100 21.700 ;
        RECT 72.500 20.000 73.100 20.700 ;
        RECT 73.600 20.000 74.710 22.000 ;
        RECT 72.800 19.970 73.050 20.000 ;
        RECT 73.630 19.970 73.880 20.000 ;
        RECT 74.460 19.970 74.710 20.000 ;
        RECT 75.290 22.000 75.540 22.075 ;
        RECT 76.120 22.000 76.370 22.075 ;
        RECT 76.950 22.000 77.200 22.075 ;
        RECT 77.780 22.000 78.030 22.075 ;
        RECT 75.290 20.000 76.400 22.000 ;
        RECT 76.900 20.000 78.030 22.000 ;
        RECT 75.290 19.970 75.540 20.000 ;
        RECT 76.120 19.970 76.370 20.000 ;
        RECT 76.950 19.970 77.200 20.000 ;
        RECT 77.780 19.970 78.030 20.000 ;
        RECT 78.610 22.000 78.860 22.075 ;
        RECT 80.170 22.000 80.420 22.075 ;
        RECT 78.610 20.000 80.420 22.000 ;
        RECT 78.610 19.970 78.860 20.000 ;
        RECT 80.170 19.970 80.420 20.000 ;
        RECT 81.000 22.000 81.250 22.075 ;
        RECT 81.830 22.000 82.080 22.075 ;
        RECT 82.660 22.000 82.910 22.075 ;
        RECT 83.490 22.000 83.740 22.075 ;
        RECT 84.320 22.000 84.570 22.075 ;
        RECT 85.150 22.000 85.400 22.075 ;
        RECT 81.000 20.000 82.200 22.000 ;
        RECT 82.660 20.000 83.800 22.000 ;
        RECT 84.300 20.000 85.400 22.000 ;
        RECT 85.980 20.200 86.230 22.075 ;
        RECT 81.000 19.970 81.250 20.000 ;
        RECT 81.830 19.970 82.080 20.000 ;
        RECT 82.660 19.970 82.910 20.000 ;
        RECT 83.490 19.970 83.740 20.000 ;
        RECT 84.320 19.970 84.570 20.000 ;
        RECT 85.150 19.970 85.400 20.000 ;
        RECT 85.900 19.800 86.300 20.200 ;
        RECT 83.800 19.400 86.300 19.800 ;
        RECT 57.640 18.765 59.240 19.210 ;
        RECT 85.850 19.000 86.550 19.100 ;
        RECT 57.640 18.310 59.140 18.765 ;
        RECT 72.850 18.500 86.550 19.000 ;
        RECT 50.340 16.795 51.840 16.810 ;
        RECT 50.320 16.510 51.840 16.795 ;
        RECT 50.320 15.610 50.550 16.510 ;
        RECT 51.610 16.505 51.840 16.510 ;
        RECT 55.140 16.010 55.370 18.310 ;
        RECT 57.720 16.010 57.950 18.310 ;
        RECT 60.140 16.010 61.140 16.310 ;
        RECT 51.040 15.910 61.140 16.010 ;
        RECT 50.990 15.610 61.140 15.910 ;
        RECT 72.950 15.900 73.350 17.900 ;
        RECT 73.880 17.800 74.130 17.890 ;
        RECT 74.710 17.800 74.960 17.890 ;
        RECT 73.880 15.900 74.960 17.800 ;
        RECT 73.050 15.785 73.300 15.900 ;
        RECT 73.880 15.785 74.130 15.900 ;
        RECT 74.710 15.785 74.960 15.900 ;
        RECT 75.540 17.800 75.790 17.890 ;
        RECT 76.370 17.800 76.620 17.890 ;
        RECT 75.540 15.900 76.620 17.800 ;
        RECT 75.540 15.785 75.790 15.900 ;
        RECT 76.370 15.785 76.620 15.900 ;
        RECT 77.200 17.800 77.450 17.890 ;
        RECT 78.030 17.800 78.280 17.890 ;
        RECT 77.200 15.900 78.280 17.800 ;
        RECT 77.200 15.785 77.450 15.900 ;
        RECT 78.030 15.785 78.280 15.900 ;
        RECT 78.860 17.300 79.110 17.890 ;
        RECT 78.860 17.200 82.700 17.300 ;
        RECT 78.860 16.100 82.750 17.200 ;
        RECT 78.860 15.785 79.110 16.100 ;
        RECT 3.700 13.385 14.260 14.000 ;
        RECT 2.090 12.865 3.050 13.095 ;
        RECT 3.700 12.800 14.200 13.385 ;
        RECT 14.890 12.865 15.850 13.095 ;
        RECT 30.140 12.710 30.370 15.210 ;
        RECT 32.720 12.710 32.950 15.210 ;
        RECT 45.160 15.110 50.550 15.610 ;
        RECT 45.160 14.710 45.390 15.110 ;
        RECT 44.140 14.235 45.390 14.710 ;
        RECT 47.590 14.310 47.990 15.110 ;
        RECT 50.320 14.510 50.550 15.110 ;
        RECT 47.740 14.235 47.970 14.310 ;
        RECT 50.320 14.235 51.340 14.510 ;
        RECT 44.140 13.910 45.240 14.235 ;
        RECT 50.440 13.990 51.340 14.235 ;
        RECT 44.150 13.760 45.110 13.910 ;
        RECT 45.440 13.760 46.400 13.990 ;
        RECT 46.730 13.760 47.690 13.990 ;
        RECT 48.020 13.760 48.980 13.990 ;
        RECT 49.310 13.760 50.270 13.990 ;
        RECT 50.440 13.810 51.560 13.990 ;
        RECT 50.600 13.760 51.560 13.810 ;
        RECT 40.480 12.980 41.100 13.440 ;
        RECT 47.580 12.980 48.200 13.440 ;
        RECT 10.150 12.100 15.150 12.400 ;
        RECT 2.650 11.200 6.250 11.600 ;
        RECT 6.450 11.400 13.650 11.800 ;
        RECT 30.140 11.210 30.440 12.710 ;
        RECT 32.720 11.495 33.040 12.710 ;
        RECT 32.740 11.210 33.040 11.495 ;
        RECT 55.140 12.310 55.370 15.610 ;
        RECT 57.720 12.310 57.950 15.610 ;
        RECT 60.140 15.310 61.140 15.610 ;
        RECT 73.050 13.600 73.300 13.735 ;
        RECT 73.880 13.600 74.130 13.735 ;
        RECT 55.140 11.310 55.440 12.310 ;
        RECT 57.720 11.495 58.040 12.310 ;
        RECT 73.050 11.700 74.130 13.600 ;
        RECT 73.050 11.630 73.300 11.700 ;
        RECT 73.880 11.630 74.130 11.700 ;
        RECT 74.710 13.600 74.960 13.735 ;
        RECT 75.540 13.600 75.790 13.735 ;
        RECT 74.710 11.700 75.790 13.600 ;
        RECT 74.710 11.630 74.960 11.700 ;
        RECT 75.540 11.630 75.790 11.700 ;
        RECT 76.370 13.600 76.620 13.735 ;
        RECT 77.200 13.600 77.450 13.735 ;
        RECT 76.370 11.700 77.450 13.600 ;
        RECT 76.370 11.630 76.620 11.700 ;
        RECT 77.200 11.630 77.450 11.700 ;
        RECT 78.030 13.600 78.280 13.735 ;
        RECT 78.860 13.600 79.110 13.735 ;
        RECT 78.030 11.700 79.110 13.600 ;
        RECT 118.800 13.200 119.900 13.500 ;
        RECT 82.150 12.700 122.150 13.200 ;
        RECT 82.200 12.600 122.150 12.700 ;
        RECT 118.800 12.400 119.900 12.600 ;
        RECT 78.030 11.630 78.280 11.700 ;
        RECT 78.860 11.630 79.110 11.700 ;
        RECT 57.740 11.310 58.040 11.495 ;
        RECT 29.140 11.205 33.940 11.210 ;
        RECT 54.040 11.205 58.940 11.310 ;
        RECT 29.130 11.010 33.960 11.205 ;
        RECT 54.040 11.010 58.960 11.205 ;
        RECT 29.130 10.975 30.090 11.010 ;
        RECT 33.000 10.975 33.960 11.010 ;
        RECT 54.130 10.975 55.090 11.010 ;
        RECT 58.000 10.975 58.960 11.010 ;
        RECT 13.450 10.400 15.050 10.800 ;
        RECT 26.840 10.510 27.840 10.710 ;
        RECT 26.840 10.110 35.590 10.510 ;
        RECT 0.800 1.050 2.400 9.850 ;
        RECT 13.350 9.800 13.850 9.900 ;
        RECT 3.000 9.600 13.850 9.800 ;
        RECT 14.410 9.700 15.700 9.750 ;
        RECT 26.840 9.710 27.840 10.110 ;
        RECT 3.010 9.520 3.970 9.600 ;
        RECT 4.910 9.520 5.870 9.600 ;
        RECT 6.810 9.520 7.770 9.600 ;
        RECT 8.710 9.520 9.670 9.600 ;
        RECT 10.610 9.520 11.570 9.600 ;
        RECT 12.510 9.520 13.470 9.600 ;
        RECT 14.300 9.500 15.700 9.700 ;
        RECT 2.730 9.350 2.960 9.360 ;
        RECT 4.020 9.350 4.250 9.360 ;
        RECT 4.630 9.350 4.860 9.360 ;
        RECT 5.920 9.350 6.150 9.360 ;
        RECT 2.650 8.450 3.050 9.350 ;
        RECT 2.730 8.360 2.960 8.450 ;
        RECT 4.020 8.360 4.860 9.350 ;
        RECT 5.850 8.450 6.250 9.350 ;
        RECT 6.530 9.250 6.760 9.360 ;
        RECT 7.820 9.350 8.050 9.360 ;
        RECT 8.430 9.350 8.660 9.360 ;
        RECT 6.450 8.450 6.850 9.250 ;
        RECT 5.920 8.360 6.150 8.450 ;
        RECT 6.530 8.360 6.760 8.450 ;
        RECT 7.820 8.360 8.660 9.350 ;
        RECT 9.720 9.300 9.950 9.360 ;
        RECT 10.330 9.350 10.560 9.360 ;
        RECT 11.620 9.350 11.850 9.360 ;
        RECT 12.230 9.350 12.460 9.360 ;
        RECT 9.550 8.400 9.950 9.300 ;
        RECT 9.720 8.360 9.950 8.400 ;
        RECT 4.050 8.350 4.850 8.360 ;
        RECT 7.900 8.350 8.600 8.360 ;
        RECT 10.150 8.350 10.650 9.350 ;
        RECT 11.620 8.450 12.460 9.350 ;
        RECT 13.520 9.250 13.750 9.360 ;
        RECT 11.620 8.360 11.850 8.450 ;
        RECT 12.230 8.360 12.460 8.450 ;
        RECT 13.350 8.350 13.750 9.250 ;
        RECT 3.010 7.970 3.970 8.200 ;
        RECT 4.910 7.970 5.870 8.200 ;
        RECT 6.810 7.970 7.770 8.200 ;
        RECT 8.710 7.970 9.670 8.200 ;
        RECT 10.610 7.970 11.570 8.200 ;
        RECT 12.510 7.970 13.470 8.200 ;
        RECT 3.300 7.660 3.800 7.970 ;
        RECT 5.100 7.660 5.600 7.970 ;
        RECT 7.000 7.660 7.500 7.970 ;
        RECT 9.000 7.660 9.500 7.970 ;
        RECT 10.900 7.660 11.400 7.970 ;
        RECT 12.700 7.660 13.200 7.970 ;
        RECT 3.010 7.430 3.970 7.660 ;
        RECT 4.910 7.430 5.870 7.660 ;
        RECT 6.810 7.430 7.770 7.660 ;
        RECT 8.710 7.430 9.670 7.660 ;
        RECT 10.610 7.430 11.570 7.660 ;
        RECT 12.510 7.430 13.470 7.660 ;
        RECT 5.100 7.400 5.600 7.430 ;
        RECT 7.000 7.400 7.500 7.430 ;
        RECT 9.000 7.400 9.500 7.430 ;
        RECT 10.900 7.400 11.400 7.430 ;
        RECT 12.700 7.400 13.200 7.430 ;
        RECT 2.730 7.250 2.960 7.270 ;
        RECT 4.020 7.250 4.250 7.270 ;
        RECT 4.630 7.250 4.860 7.270 ;
        RECT 5.920 7.250 6.150 7.270 ;
        RECT 2.650 6.250 3.050 7.250 ;
        RECT 4.020 6.270 4.860 7.250 ;
        RECT 5.850 6.350 6.250 7.250 ;
        RECT 6.530 7.150 6.760 7.270 ;
        RECT 7.820 7.250 8.050 7.270 ;
        RECT 8.430 7.250 8.660 7.270 ;
        RECT 6.450 6.350 6.850 7.150 ;
        RECT 5.920 6.270 6.150 6.350 ;
        RECT 6.530 6.270 6.760 6.350 ;
        RECT 7.820 6.270 8.660 7.250 ;
        RECT 9.720 7.200 9.950 7.270 ;
        RECT 10.330 7.250 10.560 7.270 ;
        RECT 11.620 7.250 11.850 7.270 ;
        RECT 12.230 7.250 12.460 7.270 ;
        RECT 13.520 7.250 13.750 7.270 ;
        RECT 9.550 6.300 9.950 7.200 ;
        RECT 9.720 6.270 9.950 6.300 ;
        RECT 4.050 6.250 4.850 6.270 ;
        RECT 7.900 6.250 8.600 6.270 ;
        RECT 10.250 6.250 10.750 7.250 ;
        RECT 11.620 6.350 12.460 7.250 ;
        RECT 13.450 6.350 13.850 7.250 ;
        RECT 11.620 6.270 11.850 6.350 ;
        RECT 12.230 6.270 12.460 6.350 ;
        RECT 13.520 6.270 13.750 6.350 ;
        RECT 3.010 5.880 3.970 6.110 ;
        RECT 4.910 5.880 5.870 6.110 ;
        RECT 6.810 5.880 7.770 6.110 ;
        RECT 8.710 5.880 9.670 6.110 ;
        RECT 10.610 5.880 11.570 6.110 ;
        RECT 12.510 5.880 13.470 6.110 ;
        RECT 3.300 5.570 3.800 5.880 ;
        RECT 5.100 5.570 5.600 5.880 ;
        RECT 7.000 5.570 7.500 5.880 ;
        RECT 9.000 5.570 9.500 5.880 ;
        RECT 10.900 5.570 11.400 5.880 ;
        RECT 12.700 5.570 13.200 5.880 ;
        RECT 3.010 5.340 3.970 5.570 ;
        RECT 4.910 5.340 5.870 5.570 ;
        RECT 6.810 5.340 7.770 5.570 ;
        RECT 8.710 5.340 9.670 5.570 ;
        RECT 10.610 5.340 11.570 5.570 ;
        RECT 12.510 5.340 13.470 5.570 ;
        RECT 2.730 5.150 2.960 5.180 ;
        RECT 4.020 5.150 4.250 5.180 ;
        RECT 4.630 5.150 4.860 5.180 ;
        RECT 5.920 5.150 6.150 5.180 ;
        RECT 2.650 4.250 3.050 5.150 ;
        RECT 2.730 4.180 2.960 4.250 ;
        RECT 4.020 4.180 4.860 5.150 ;
        RECT 5.850 4.250 6.250 5.150 ;
        RECT 6.530 5.050 6.760 5.180 ;
        RECT 7.820 5.150 8.050 5.180 ;
        RECT 8.430 5.150 8.660 5.180 ;
        RECT 6.450 4.250 6.850 5.050 ;
        RECT 5.920 4.180 6.150 4.250 ;
        RECT 6.530 4.180 6.760 4.250 ;
        RECT 7.820 4.180 8.660 5.150 ;
        RECT 9.720 5.100 9.950 5.180 ;
        RECT 10.330 5.150 10.560 5.180 ;
        RECT 11.620 5.150 11.850 5.180 ;
        RECT 12.230 5.150 12.460 5.180 ;
        RECT 13.520 5.150 13.750 5.180 ;
        RECT 9.550 4.200 9.950 5.100 ;
        RECT 10.250 4.250 10.650 5.150 ;
        RECT 11.620 4.250 12.460 5.150 ;
        RECT 13.450 4.250 13.850 5.150 ;
        RECT 9.720 4.180 9.950 4.200 ;
        RECT 10.330 4.180 10.560 4.250 ;
        RECT 11.620 4.180 11.850 4.250 ;
        RECT 12.230 4.180 12.460 4.250 ;
        RECT 13.520 4.180 13.750 4.250 ;
        RECT 4.050 4.150 4.850 4.180 ;
        RECT 7.900 4.150 8.600 4.180 ;
        RECT 3.010 3.790 3.970 4.020 ;
        RECT 4.910 3.790 5.870 4.020 ;
        RECT 6.810 3.790 7.770 4.020 ;
        RECT 8.710 3.790 9.670 4.020 ;
        RECT 10.610 3.790 11.570 4.020 ;
        RECT 12.510 3.790 13.470 4.020 ;
        RECT 3.300 3.480 3.800 3.790 ;
        RECT 5.100 3.480 5.600 3.790 ;
        RECT 7.000 3.480 7.500 3.790 ;
        RECT 9.000 3.480 9.500 3.790 ;
        RECT 10.900 3.480 11.400 3.790 ;
        RECT 12.700 3.480 13.200 3.790 ;
        RECT 3.010 3.250 3.970 3.480 ;
        RECT 4.910 3.250 5.870 3.480 ;
        RECT 6.810 3.250 7.770 3.480 ;
        RECT 8.710 3.250 9.670 3.480 ;
        RECT 10.610 3.250 11.570 3.480 ;
        RECT 12.510 3.250 13.470 3.480 ;
        RECT 2.730 3.050 2.960 3.090 ;
        RECT 4.020 3.050 4.250 3.090 ;
        RECT 4.630 3.050 4.860 3.090 ;
        RECT 5.920 3.050 6.150 3.090 ;
        RECT 2.650 2.150 3.050 3.050 ;
        RECT 4.020 2.150 4.860 3.050 ;
        RECT 5.850 2.150 6.250 3.050 ;
        RECT 6.530 2.950 6.760 3.090 ;
        RECT 7.820 3.050 8.050 3.090 ;
        RECT 8.430 3.050 8.660 3.090 ;
        RECT 6.450 2.150 6.850 2.950 ;
        RECT 2.730 2.090 2.960 2.150 ;
        RECT 4.020 2.090 4.250 2.150 ;
        RECT 4.630 2.090 4.860 2.150 ;
        RECT 5.920 2.090 6.150 2.150 ;
        RECT 6.530 2.090 6.760 2.150 ;
        RECT 7.820 2.090 8.660 3.050 ;
        RECT 9.720 3.000 9.950 3.090 ;
        RECT 10.330 3.050 10.560 3.090 ;
        RECT 11.620 3.050 11.850 3.090 ;
        RECT 12.230 3.050 12.460 3.090 ;
        RECT 13.520 3.050 13.750 3.090 ;
        RECT 9.550 2.100 9.950 3.000 ;
        RECT 10.250 2.150 10.650 3.050 ;
        RECT 11.620 2.150 12.460 3.050 ;
        RECT 13.450 2.150 13.850 3.050 ;
        RECT 9.720 2.090 9.950 2.100 ;
        RECT 10.330 2.090 10.560 2.150 ;
        RECT 11.620 2.090 11.850 2.150 ;
        RECT 12.230 2.090 12.460 2.150 ;
        RECT 13.520 2.090 13.750 2.150 ;
        RECT 7.900 2.050 8.600 2.090 ;
        RECT 3.010 1.700 3.970 1.930 ;
        RECT 4.910 1.700 5.870 1.930 ;
        RECT 6.810 1.700 7.770 1.930 ;
        RECT 8.710 1.700 9.670 1.930 ;
        RECT 10.610 1.700 11.570 1.930 ;
        RECT 12.510 1.700 13.470 1.930 ;
        RECT 5.440 1.050 6.660 1.230 ;
        RECT 10.040 1.050 11.260 1.230 ;
        RECT 14.100 1.050 15.700 9.500 ;
        RECT 85.850 9.200 86.250 9.300 ;
        RECT 26.840 9.100 27.840 9.110 ;
        RECT 24.900 8.910 27.840 9.100 ;
        RECT 85.850 9.000 86.300 9.200 ;
        RECT 85.980 8.970 86.270 9.000 ;
        RECT 24.900 8.310 39.990 8.910 ;
        RECT 69.930 8.550 72.500 8.900 ;
        RECT 85.350 8.765 85.900 8.800 ;
        RECT 24.900 8.110 27.840 8.310 ;
        RECT 24.900 8.100 27.800 8.110 ;
        RECT 69.930 8.000 84.900 8.550 ;
        RECT 69.930 7.900 72.500 8.000 ;
        RECT 71.500 7.800 72.500 7.900 ;
        RECT 71.500 7.000 72.500 7.300 ;
        RECT 71.500 6.520 83.570 7.000 ;
        RECT 71.500 6.500 73.200 6.520 ;
        RECT 71.500 6.300 72.600 6.500 ;
        RECT 72.100 6.100 72.600 6.300 ;
        RECT 73.945 5.980 74.235 6.025 ;
        RECT 75.835 5.980 76.125 6.025 ;
        RECT 78.955 5.980 79.245 6.025 ;
        RECT 73.945 5.840 79.245 5.980 ;
        RECT 85.350 5.900 86.020 8.765 ;
        RECT 73.945 5.795 74.235 5.840 ;
        RECT 75.835 5.795 76.125 5.840 ;
        RECT 78.955 5.795 79.245 5.840 ;
        RECT 85.790 5.765 86.020 5.900 ;
        RECT 86.230 8.700 86.460 8.765 ;
        RECT 86.770 8.700 87.030 8.760 ;
        RECT 86.230 8.600 87.200 8.700 ;
        RECT 86.230 8.200 87.250 8.600 ;
        RECT 86.230 8.000 87.200 8.200 ;
        RECT 86.230 7.600 87.250 8.000 ;
        RECT 86.230 7.300 87.200 7.600 ;
        RECT 86.230 6.900 87.250 7.300 ;
        RECT 86.230 6.600 87.200 6.900 ;
        RECT 86.230 6.200 87.250 6.600 ;
        RECT 86.230 5.900 87.200 6.200 ;
        RECT 86.230 5.765 86.460 5.900 ;
        RECT 86.770 5.840 87.030 5.900 ;
        RECT 65.400 5.500 72.500 5.600 ;
        RECT 85.980 5.500 86.270 5.560 ;
        RECT 65.350 5.400 72.500 5.500 ;
        RECT 73.070 5.400 73.330 5.460 ;
        RECT 65.350 5.100 73.330 5.400 ;
        RECT 73.540 5.300 73.830 5.345 ;
        RECT 75.375 5.300 75.665 5.345 ;
        RECT 78.955 5.300 79.245 5.345 ;
        RECT 73.540 5.160 79.245 5.300 ;
        RECT 73.540 5.115 73.830 5.160 ;
        RECT 75.375 5.115 75.665 5.160 ;
        RECT 78.955 5.115 79.245 5.160 ;
        RECT 65.350 4.600 72.500 5.100 ;
        RECT 73.070 5.040 73.330 5.100 ;
        RECT 80.035 5.005 80.325 5.320 ;
        RECT 83.190 5.300 83.510 5.330 ;
        RECT 84.450 5.300 84.950 5.400 ;
        RECT 85.900 5.300 86.350 5.500 ;
        RECT 83.190 5.100 84.950 5.300 ;
        RECT 85.950 5.200 86.350 5.300 ;
        RECT 83.190 5.070 83.510 5.100 ;
        RECT 76.735 5.000 77.385 5.005 ;
        RECT 74.400 4.650 74.900 5.000 ;
        RECT 76.650 4.960 77.385 5.000 ;
        RECT 80.035 4.960 80.625 5.005 ;
        RECT 84.450 5.000 84.950 5.100 ;
        RECT 76.650 4.820 80.625 4.960 ;
        RECT 76.650 4.775 77.385 4.820 ;
        RECT 80.335 4.775 80.625 4.820 ;
        RECT 81.640 4.800 82.060 4.830 ;
        RECT 76.650 4.700 77.050 4.775 ;
        RECT 81.640 4.500 84.350 4.800 ;
        RECT 81.640 4.470 82.060 4.500 ;
        RECT 72.990 3.800 83.570 4.280 ;
        RECT 85.950 3.800 86.350 3.900 ;
        RECT 85.900 3.600 86.350 3.800 ;
        RECT 74.450 3.300 85.650 3.600 ;
        RECT 85.980 3.530 86.270 3.600 ;
        RECT 85.790 3.300 86.020 3.370 ;
        RECT 85.250 3.250 86.020 3.300 ;
        RECT 71.500 2.500 72.500 2.800 ;
        RECT 71.500 2.200 77.050 2.500 ;
        RECT 85.350 2.400 86.020 3.250 ;
        RECT 85.790 2.370 86.020 2.400 ;
        RECT 86.230 3.300 86.460 3.370 ;
        RECT 86.230 2.400 87.300 3.300 ;
        RECT 86.230 2.370 86.460 2.400 ;
        RECT 86.700 2.300 87.300 2.400 ;
        RECT 85.980 2.200 86.270 2.210 ;
        RECT 71.500 1.800 72.500 2.200 ;
        RECT 85.900 2.000 86.300 2.200 ;
        RECT 85.980 1.980 86.270 2.000 ;
        RECT 0.800 0.000 15.700 1.050 ;
        RECT 78.600 0.800 79.600 1.000 ;
        RECT 72.900 0.700 87.100 0.800 ;
        RECT 72.900 0.100 87.150 0.700 ;
        RECT 72.900 0.000 87.100 0.100 ;
        RECT 80.150 -0.100 80.950 0.000 ;
        RECT 0.290 -8.780 80.490 -7.980 ;
        RECT 0.690 -9.780 80.490 -8.780 ;
        RECT 0.290 -10.180 80.490 -9.780 ;
        RECT 24.790 -10.800 25.790 -10.780 ;
        RECT 21.790 -10.980 22.790 -10.880 ;
        RECT 21.740 -11.480 22.840 -10.980 ;
        RECT 21.800 -11.900 22.800 -11.480 ;
        RECT 24.750 -11.500 25.850 -10.800 ;
        RECT 24.790 -11.880 25.790 -11.500 ;
        RECT 65.390 -11.880 66.390 -10.780 ;
        RECT 68.490 -11.880 69.290 -10.880 ;
        RECT 70.040 -11.480 70.940 -10.880 ;
        RECT 70.090 -11.880 70.890 -11.480 ;
        RECT 71.490 -11.880 72.490 -10.780 ;
      LAYER via ;
        RECT 34.700 34.400 36.300 35.800 ;
        RECT 1.600 26.500 2.000 27.000 ;
        RECT 8.000 26.500 8.600 27.000 ;
        RECT 17.500 26.600 20.000 27.400 ;
        RECT 31.440 27.210 31.740 27.810 ;
        RECT 40.940 27.210 41.440 27.710 ;
        RECT 43.800 27.700 44.800 29.500 ;
        RECT 46.640 27.210 47.140 27.710 ;
        RECT 56.340 27.110 56.640 27.610 ;
        RECT 20.200 26.500 20.700 27.000 ;
        RECT 8.000 24.200 8.600 24.800 ;
        RECT 11.800 22.900 12.200 24.000 ;
        RECT 20.200 24.200 20.700 24.800 ;
        RECT 16.400 23.100 16.900 23.700 ;
        RECT 13.100 22.400 13.600 22.700 ;
        RECT 1.600 21.100 2.000 21.500 ;
        RECT 11.800 21.000 12.200 21.500 ;
        RECT 14.600 20.900 15.100 21.400 ;
        RECT 4.200 19.000 4.700 19.300 ;
        RECT 13.100 19.000 13.600 19.300 ;
        RECT 31.340 24.410 31.840 25.610 ;
        RECT 40.940 26.010 41.440 26.410 ;
        RECT 42.340 25.410 42.740 25.910 ;
        RECT 45.540 25.810 45.940 26.210 ;
        RECT 46.740 25.410 47.140 26.010 ;
        RECT 43.840 23.710 44.240 24.110 ;
        RECT 52.640 23.710 53.040 24.110 ;
        RECT 43.840 23.210 44.240 23.510 ;
        RECT 42.340 22.610 42.740 23.010 ;
        RECT 45.540 22.610 45.940 23.010 ;
        RECT 44.040 21.610 44.340 22.010 ;
        RECT 45.540 21.110 45.840 21.410 ;
        RECT 35.240 20.510 35.540 20.810 ;
        RECT 45.540 20.510 45.840 20.810 ;
        RECT 41.940 20.010 42.340 20.310 ;
        RECT 44.040 20.010 44.340 20.310 ;
        RECT 13.100 17.100 13.600 17.700 ;
        RECT 39.540 18.710 39.940 19.110 ;
        RECT 40.540 18.510 41.040 19.010 ;
        RECT 41.940 18.810 42.240 19.310 ;
        RECT 56.340 23.410 56.640 26.210 ;
        RECT 44.340 18.110 44.640 18.410 ;
        RECT 45.740 18.110 46.040 19.010 ;
        RECT 50.940 17.510 51.240 17.810 ;
        RECT 16.400 14.700 17.000 15.200 ;
        RECT 21.900 14.500 22.800 15.500 ;
        RECT 26.900 14.600 27.700 15.400 ;
        RECT 44.340 15.310 44.640 15.610 ;
        RECT 60.200 26.200 61.000 27.000 ;
        RECT 68.600 26.200 69.200 27.000 ;
        RECT 71.500 26.200 72.200 27.000 ;
        RECT 86.600 28.500 87.500 29.400 ;
        RECT 86.800 27.200 87.300 27.600 ;
        RECT 71.600 20.800 72.300 21.600 ;
        RECT 79.300 20.100 79.700 21.900 ;
        RECT 83.900 19.400 84.300 19.700 ;
        RECT 72.900 18.500 73.400 19.000 ;
        RECT 79.300 18.600 79.700 19.000 ;
        RECT 85.900 18.500 86.500 19.100 ;
        RECT 51.040 15.610 51.340 15.910 ;
        RECT 52.640 15.710 52.940 16.010 ;
        RECT 13.100 12.900 13.500 13.900 ;
        RECT 47.640 14.310 47.940 15.510 ;
        RECT 40.540 13.010 41.040 13.410 ;
        RECT 47.640 13.010 48.140 13.410 ;
        RECT 10.200 12.100 10.500 12.400 ;
        RECT 14.600 12.100 15.100 12.400 ;
        RECT 2.700 11.200 3.000 11.600 ;
        RECT 4.200 11.200 4.700 11.500 ;
        RECT 5.900 11.200 6.200 11.600 ;
        RECT 6.500 11.400 6.800 11.800 ;
        RECT 9.700 11.400 10.000 11.800 ;
        RECT 13.100 11.400 13.600 11.800 ;
        RECT 60.200 15.400 61.000 16.200 ;
        RECT 73.000 15.900 73.300 17.900 ;
        RECT 82.200 16.100 82.700 17.200 ;
        RECT 82.200 12.700 82.800 13.200 ;
        RECT 85.900 12.600 86.300 13.200 ;
        RECT 118.900 12.500 119.800 13.400 ;
        RECT 13.500 10.400 13.800 10.800 ;
        RECT 14.600 10.400 15.000 10.800 ;
        RECT 13.400 9.600 13.800 9.900 ;
        RECT 26.900 9.800 27.700 10.600 ;
        RECT 35.240 10.110 35.540 10.510 ;
        RECT 2.700 8.450 3.000 9.350 ;
        RECT 4.100 8.350 4.800 9.350 ;
        RECT 5.900 8.450 6.200 9.350 ;
        RECT 6.500 8.450 6.800 9.250 ;
        RECT 7.900 8.450 8.400 9.150 ;
        RECT 9.600 8.400 9.900 9.300 ;
        RECT 10.200 8.350 10.600 9.350 ;
        RECT 11.700 8.450 12.300 9.250 ;
        RECT 13.400 8.350 13.700 9.250 ;
        RECT 2.700 6.250 3.000 7.250 ;
        RECT 4.100 6.250 4.800 7.250 ;
        RECT 5.900 6.350 6.200 7.250 ;
        RECT 6.500 6.350 6.800 7.150 ;
        RECT 8.000 6.350 8.500 7.050 ;
        RECT 9.600 6.300 9.900 7.200 ;
        RECT 10.300 6.250 10.700 7.250 ;
        RECT 11.700 6.350 12.300 7.150 ;
        RECT 13.500 6.350 13.800 7.250 ;
        RECT 2.700 4.250 3.000 5.150 ;
        RECT 4.100 4.150 4.800 5.150 ;
        RECT 5.900 4.250 6.200 5.150 ;
        RECT 6.500 4.250 6.800 5.050 ;
        RECT 8.000 4.250 8.500 4.950 ;
        RECT 9.600 4.200 9.900 5.100 ;
        RECT 10.300 4.250 10.600 5.150 ;
        RECT 11.700 4.250 12.300 5.050 ;
        RECT 13.500 4.250 13.800 5.150 ;
        RECT 2.700 2.150 3.000 3.050 ;
        RECT 4.100 2.150 4.800 3.050 ;
        RECT 5.900 2.150 6.200 3.050 ;
        RECT 6.500 2.150 6.800 2.950 ;
        RECT 8.000 2.150 8.500 2.850 ;
        RECT 9.600 2.100 9.900 3.000 ;
        RECT 10.300 2.150 10.600 3.050 ;
        RECT 11.700 2.150 12.300 2.950 ;
        RECT 13.500 2.150 13.800 3.050 ;
        RECT 85.900 9.000 86.200 9.300 ;
        RECT 25.000 8.200 25.600 9.000 ;
        RECT 39.540 8.310 39.940 8.910 ;
        RECT 70.100 7.900 70.800 8.900 ;
        RECT 84.500 8.000 84.850 8.550 ;
        RECT 71.700 6.400 72.300 7.100 ;
        RECT 85.400 5.900 85.700 8.800 ;
        RECT 86.800 8.200 87.200 8.600 ;
        RECT 86.800 7.600 87.200 8.000 ;
        RECT 86.800 6.900 87.200 7.300 ;
        RECT 86.800 6.200 87.200 6.600 ;
        RECT 65.400 4.600 66.300 5.500 ;
        RECT 74.450 4.650 74.850 5.000 ;
        RECT 76.700 4.700 77.000 5.000 ;
        RECT 84.500 5.000 84.900 5.400 ;
        RECT 86.000 5.200 86.300 5.500 ;
        RECT 83.900 4.500 84.300 4.800 ;
        RECT 73.100 3.800 73.500 4.200 ;
        RECT 86.000 3.600 86.300 3.900 ;
        RECT 74.500 3.300 74.800 3.600 ;
        RECT 85.300 3.250 85.600 3.550 ;
        RECT 71.700 1.800 72.300 2.700 ;
        RECT 76.700 2.200 77.000 2.500 ;
        RECT 86.600 2.400 87.100 3.100 ;
        RECT 1.000 0.200 2.400 0.800 ;
        RECT 4.200 0.450 4.700 0.950 ;
        RECT 7.900 0.350 8.500 1.050 ;
        RECT 11.700 0.350 12.400 1.050 ;
        RECT 73.000 0.100 73.500 0.800 ;
        RECT 78.200 0.100 79.500 0.700 ;
        RECT 86.600 0.100 87.100 0.700 ;
        RECT 0.990 -9.580 2.290 -8.080 ;
        RECT 40.640 -8.590 40.940 -8.290 ;
        RECT 47.740 -8.590 48.040 -8.290 ;
        RECT 78.390 -9.380 79.390 -8.180 ;
        RECT 21.790 -11.480 22.790 -10.980 ;
        RECT 24.800 -11.500 25.800 -10.800 ;
        RECT 65.490 -11.380 66.290 -10.880 ;
        RECT 68.590 -11.380 69.190 -10.980 ;
        RECT 70.090 -11.480 70.890 -10.880 ;
        RECT 71.590 -11.380 72.390 -10.880 ;
      LAYER met2 ;
        RECT 34.700 34.350 36.300 35.850 ;
        RECT 31.440 27.810 31.740 27.860 ;
        RECT 1.600 21.050 2.000 27.050 ;
        RECT 8.000 24.150 8.600 27.050 ;
        RECT 17.500 26.550 20.000 27.450 ;
        RECT 20.200 24.150 20.700 27.050 ;
        RECT 31.340 24.360 31.840 27.810 ;
        RECT 40.940 25.960 41.440 27.760 ;
        RECT 43.800 27.650 44.800 29.550 ;
        RECT 86.600 28.450 87.500 29.450 ;
        RECT 11.800 20.950 12.200 24.050 ;
        RECT 2.700 2.050 3.000 11.650 ;
        RECT 4.200 11.150 4.700 19.350 ;
        RECT 0.800 -6.920 2.500 0.900 ;
        RECT 4.100 0.350 4.800 9.400 ;
        RECT 5.900 2.050 6.200 11.650 ;
        RECT 6.500 2.050 6.800 11.850 ;
        RECT 9.700 9.350 10.000 11.850 ;
        RECT 7.900 0.300 8.500 9.250 ;
        RECT 9.600 8.350 10.000 9.350 ;
        RECT 9.700 7.250 10.000 8.350 ;
        RECT 9.600 6.250 10.000 7.250 ;
        RECT 9.700 5.150 10.000 6.250 ;
        RECT 9.600 4.150 10.000 5.150 ;
        RECT 9.700 3.050 10.000 4.150 ;
        RECT 9.600 2.050 10.000 3.050 ;
        RECT 10.200 9.400 10.500 12.450 ;
        RECT 13.100 11.350 13.600 22.750 ;
        RECT 14.600 11.950 15.100 21.450 ;
        RECT 16.400 14.650 17.000 23.800 ;
        RECT 42.340 22.560 42.740 26.010 ;
        RECT 43.840 23.160 44.240 24.160 ;
        RECT 45.540 22.560 45.940 26.260 ;
        RECT 46.640 25.410 47.140 27.760 ;
        RECT 46.740 25.360 47.140 25.410 ;
        RECT 13.500 9.950 13.800 10.850 ;
        RECT 14.600 10.350 15.000 11.950 ;
        RECT 13.400 9.550 13.800 9.950 ;
        RECT 10.200 8.300 10.600 9.400 ;
        RECT 10.200 7.300 10.500 8.300 ;
        RECT 10.200 6.200 10.700 7.300 ;
        RECT 10.200 5.200 10.500 6.200 ;
        RECT 10.200 4.200 10.600 5.200 ;
        RECT 10.200 3.100 10.500 4.200 ;
        RECT 10.200 2.100 10.600 3.100 ;
        RECT 10.200 1.750 10.500 2.100 ;
        RECT 11.700 0.300 12.400 9.350 ;
        RECT 13.500 9.300 13.800 9.550 ;
        RECT 13.400 8.300 13.800 9.300 ;
        RECT 13.500 1.850 13.800 8.300 ;
        RECT 21.800 -6.920 22.800 15.670 ;
        RECT 26.800 9.700 27.800 15.500 ;
        RECT 35.240 10.060 35.540 20.860 ;
        RECT 0.790 -8.670 2.500 -6.920 ;
        RECT 21.790 -8.170 22.800 -6.920 ;
        RECT 0.790 -9.780 2.490 -8.670 ;
        RECT 21.790 -11.530 22.790 -8.170 ;
        RECT 24.900 -10.750 25.700 9.100 ;
        RECT 39.540 8.260 39.940 19.160 ;
        RECT 40.540 -8.690 41.040 19.060 ;
        RECT 41.940 18.810 42.340 20.360 ;
        RECT 44.040 19.960 44.340 22.060 ;
        RECT 45.540 21.310 45.840 21.460 ;
        RECT 45.540 20.410 45.940 21.310 ;
        RECT 45.740 19.010 46.040 19.060 ;
        RECT 41.940 18.760 42.240 18.810 ;
        RECT 44.240 15.210 44.740 18.510 ;
        RECT 45.640 11.360 46.140 19.010 ;
        RECT 50.940 17.810 51.240 17.860 ;
        RECT 50.940 15.610 51.340 17.810 ;
        RECT 45.040 9.860 47.140 11.360 ;
        RECT 47.640 -8.690 48.140 15.610 ;
        RECT 51.040 15.560 51.340 15.610 ;
        RECT 52.640 10.410 53.040 24.160 ;
        RECT 56.240 23.210 56.740 27.710 ;
        RECT 86.800 27.600 87.300 27.650 ;
        RECT 60.100 15.300 61.100 27.100 ;
        RECT 51.640 8.910 54.040 10.410 ;
        RECT 65.400 -6.920 66.400 5.600 ;
        RECT 68.500 -6.920 69.300 27.100 ;
        RECT 71.400 20.700 72.300 27.100 ;
        RECT 72.900 15.800 73.400 19.050 ;
        RECT 79.300 18.400 79.800 22.000 ;
        RECT 82.200 12.600 82.800 17.400 ;
        RECT 70.100 8.900 70.800 8.950 ;
        RECT 70.100 -6.920 70.900 8.900 ;
        RECT 71.500 -6.920 72.500 7.300 ;
        RECT 74.450 4.600 74.850 5.050 ;
        RECT 73.100 4.200 73.500 4.250 ;
        RECT 73.000 0.050 73.500 4.200 ;
        RECT 74.500 3.650 74.700 4.600 ;
        RECT 74.500 3.250 74.800 3.650 ;
        RECT 76.700 2.150 77.000 5.050 ;
        RECT 83.900 4.450 84.300 19.750 ;
        RECT 85.900 18.450 86.500 19.150 ;
        RECT 85.900 9.000 86.300 13.250 ;
        RECT 85.900 8.950 86.200 9.000 ;
        RECT 84.500 5.450 84.850 8.600 ;
        RECT 84.500 4.950 84.900 5.450 ;
        RECT 85.400 3.600 85.700 8.850 ;
        RECT 86.700 5.900 87.300 27.600 ;
        RECT 118.800 12.400 119.900 13.500 ;
        RECT 85.300 3.200 85.700 3.600 ;
        RECT 86.000 3.550 86.300 5.550 ;
        RECT 85.400 2.400 85.700 3.200 ;
        RECT 78.000 -6.920 79.700 1.000 ;
        RECT 86.600 0.050 87.100 4.000 ;
        RECT 65.390 -8.100 66.400 -6.920 ;
        RECT 68.490 -8.100 69.300 -6.920 ;
        RECT 70.090 -8.100 70.900 -6.920 ;
        RECT 71.490 -8.100 72.500 -6.920 ;
        RECT 24.800 -11.550 25.800 -10.750 ;
        RECT 65.390 -11.480 66.390 -8.100 ;
        RECT 68.490 -11.480 69.290 -8.100 ;
        RECT 70.090 -11.530 70.890 -8.100 ;
        RECT 71.490 -11.480 72.490 -8.100 ;
        RECT 77.990 -8.150 79.700 -6.920 ;
        RECT 77.990 -9.780 79.690 -8.150 ;
      LAYER via2 ;
        RECT 34.700 34.400 36.300 35.800 ;
        RECT 17.500 26.600 20.000 27.400 ;
        RECT 43.800 27.700 44.800 29.500 ;
        RECT 86.600 28.500 87.500 29.400 ;
        RECT 45.040 9.910 47.140 11.310 ;
        RECT 51.740 9.010 53.940 10.310 ;
        RECT 85.900 18.500 86.500 19.100 ;
        RECT 118.900 12.500 119.800 13.400 ;
        RECT 86.600 0.200 87.100 0.700 ;
      LAYER met3 ;
        RECT 34.650 34.375 36.350 35.825 ;
        RECT 34.900 28.500 87.600 29.700 ;
        RECT 43.600 27.700 45.000 28.500 ;
        RECT 86.550 28.475 87.550 28.500 ;
        RECT 43.750 27.675 44.850 27.700 ;
        RECT 17.450 27.400 20.050 27.425 ;
        RECT 17.400 26.500 36.250 27.400 ;
        RECT 17.400 26.400 36.100 26.500 ;
        RECT 85.800 18.400 86.600 19.200 ;
        RECT 45.040 11.335 47.140 11.410 ;
        RECT 44.990 9.885 47.190 11.335 ;
        RECT 45.040 7.510 47.140 9.885 ;
        RECT 51.640 8.910 54.040 10.410 ;
        RECT 26.840 -7.890 58.700 7.510 ;
        RECT 88.600 0.800 116.200 29.260 ;
        RECT 118.800 12.400 119.900 13.500 ;
        RECT 120.500 0.800 148.100 29.260 ;
        RECT 86.400 0.200 148.100 0.800 ;
        RECT 86.400 0.000 122.900 0.200 ;
      LAYER via3 ;
        RECT 34.700 34.400 36.300 35.800 ;
        RECT 35.000 28.600 36.300 29.600 ;
        RECT 34.600 26.500 36.200 27.400 ;
        RECT 85.900 18.500 86.500 19.100 ;
        RECT 51.740 9.010 53.940 10.310 ;
        RECT 58.280 -7.750 58.600 7.370 ;
        RECT 118.900 12.500 119.800 13.400 ;
        RECT 88.740 0.300 116.060 0.620 ;
        RECT 120.640 0.300 147.960 0.620 ;
      LAYER met4 ;
        RECT 34.500 32.005 36.400 36.200 ;
        RECT 34.495 31.395 36.400 32.005 ;
        RECT 34.500 25.750 36.400 31.395 ;
        RECT 88.995 19.200 115.805 28.865 ;
        RECT 84.700 17.000 115.805 19.200 ;
        RECT 51.640 8.910 54.040 10.410 ;
        RECT 51.740 7.115 53.940 8.910 ;
        RECT 27.235 -7.495 56.845 7.115 ;
        RECT 58.200 -7.830 58.680 7.450 ;
        RECT 88.995 2.055 115.805 17.000 ;
        RECT 120.895 14.000 147.705 28.865 ;
        RECT 119.600 13.500 147.705 14.000 ;
        RECT 118.800 12.400 147.705 13.500 ;
        RECT 119.600 11.800 147.705 12.400 ;
        RECT 120.895 2.055 147.705 11.800 ;
        RECT 88.660 0.220 116.140 0.700 ;
        RECT 120.560 0.220 148.040 0.700 ;
  END
END device_without_rf
END LIBRARY

