magic
tech sky130A
magscale 1 2
timestamp 1657057508
<< nwell >>
rect -554 -419 554 419
<< pmos >>
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
<< pdiff >>
rect -416 188 -358 200
rect -416 -188 -404 188
rect -370 -188 -358 188
rect -416 -200 -358 -188
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
rect 358 188 416 200
rect 358 -188 370 188
rect 404 -188 416 188
rect 358 -200 416 -188
<< pdiffc >>
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
<< nsubdiff >>
rect -518 349 -422 383
rect 422 349 518 383
rect -518 287 -484 349
rect 484 287 518 349
rect -518 -349 -484 -287
rect 484 -349 518 -287
rect -518 -383 -422 -349
rect 422 -383 518 -349
<< nsubdiffcont >>
rect -422 349 422 383
rect -518 -287 -484 287
rect 484 -287 518 287
rect -422 -383 422 -349
<< poly >>
rect -358 281 -158 297
rect -358 247 -342 281
rect -174 247 -158 281
rect -358 200 -158 247
rect -100 281 100 297
rect -100 247 -84 281
rect 84 247 100 281
rect -100 200 100 247
rect 158 281 358 297
rect 158 247 174 281
rect 342 247 358 281
rect 158 200 358 247
rect -358 -247 -158 -200
rect -358 -281 -342 -247
rect -174 -281 -158 -247
rect -358 -297 -158 -281
rect -100 -247 100 -200
rect -100 -281 -84 -247
rect 84 -281 100 -247
rect -100 -297 100 -281
rect 158 -247 358 -200
rect 158 -281 174 -247
rect 342 -281 358 -247
rect 158 -297 358 -281
<< polycont >>
rect -342 247 -174 281
rect -84 247 84 281
rect 174 247 342 281
rect -342 -281 -174 -247
rect -84 -281 84 -247
rect 174 -281 342 -247
<< locali >>
rect -518 287 -484 383
rect 484 287 518 383
rect -358 247 -342 281
rect -174 247 -158 281
rect -100 247 -84 281
rect 84 247 100 281
rect 158 247 174 281
rect 342 247 358 281
rect -404 188 -370 204
rect -404 -204 -370 -188
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect 370 188 404 204
rect 370 -204 404 -188
rect -358 -281 -342 -247
rect -174 -281 -158 -247
rect -100 -281 -84 -247
rect 84 -281 100 -247
rect 158 -281 174 -247
rect 342 -281 358 -247
rect -518 -349 -484 -287
rect 484 -349 518 -287
rect -518 -383 -422 -349
rect 422 -383 518 -349
<< viali >>
rect -484 349 -422 383
rect -422 349 422 383
rect 422 349 484 383
rect -342 247 -174 281
rect -84 247 84 281
rect 174 247 342 281
rect -404 21 -370 171
rect -146 -75 -112 75
rect 112 21 146 171
rect 370 -75 404 75
rect -342 -281 -174 -247
rect -84 -281 84 -247
rect 174 -281 342 -247
<< metal1 >>
rect -496 383 496 389
rect -496 349 -484 383
rect 484 349 496 383
rect -496 343 496 349
rect -354 281 -162 287
rect -354 247 -342 281
rect -174 247 -162 281
rect -354 241 -162 247
rect -96 281 96 287
rect -96 247 -84 281
rect 84 247 96 281
rect -96 241 96 247
rect 162 281 354 287
rect 162 247 174 281
rect 342 247 354 281
rect 162 241 354 247
rect -410 171 -364 183
rect -410 21 -404 171
rect -370 21 -364 171
rect 106 171 152 183
rect -410 9 -364 21
rect -152 75 -106 87
rect -152 -75 -146 75
rect -112 -75 -106 75
rect 106 21 112 171
rect 146 21 152 171
rect 106 9 152 21
rect 364 75 410 87
rect -152 -87 -106 -75
rect 364 -75 370 75
rect 404 -75 410 75
rect 364 -87 410 -75
rect -354 -247 -162 -241
rect -354 -281 -342 -247
rect -174 -281 -162 -247
rect -354 -287 -162 -281
rect -96 -247 96 -241
rect -96 -281 -84 -247
rect 84 -281 96 -247
rect -96 -287 96 -281
rect 162 -247 354 -241
rect 162 -281 174 -247
rect 342 -281 354 -247
rect 162 -287 354 -281
<< properties >>
string FIXED_BBOX -501 -366 501 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
