magic
tech sky130A
magscale 1 2
timestamp 1657129226
<< nwell >>
rect 3200 3900 3792 4738
rect 8020 3900 8612 4738
rect 2500 2780 3092 3618
rect 4700 3020 4800 3180
rect 3020 1660 3612 2498
rect 4460 1880 4472 2180
rect 6400 1660 6992 2498
<< pwell >>
rect 11000 1480 11592 5026
<< nmos >>
rect 11196 4616 11396 4816
rect 11196 4198 11396 4398
rect 11196 3780 11396 3980
rect 11196 3362 11396 3562
rect 11196 2944 11396 3144
rect 11196 2526 11396 2726
rect 11196 2108 11396 2308
rect 11196 1690 11396 1890
<< pmos >>
rect 3396 4119 3596 4519
rect 8216 4119 8416 4519
rect 2696 2999 2896 3399
rect 4700 3020 4800 3180
rect 3216 1879 3416 2279
rect 6596 1879 6796 2279
<< ndiff >>
rect 11138 4804 11196 4816
rect 11138 4628 11150 4804
rect 11184 4628 11196 4804
rect 11138 4616 11196 4628
rect 11396 4804 11454 4816
rect 11396 4628 11408 4804
rect 11442 4628 11454 4804
rect 11396 4616 11454 4628
rect 11138 4386 11196 4398
rect 11138 4210 11150 4386
rect 11184 4210 11196 4386
rect 11138 4198 11196 4210
rect 11396 4386 11454 4398
rect 11396 4210 11408 4386
rect 11442 4210 11454 4386
rect 11396 4198 11454 4210
rect 11138 3968 11196 3980
rect 11138 3792 11150 3968
rect 11184 3792 11196 3968
rect 11138 3780 11196 3792
rect 11396 3968 11454 3980
rect 11396 3792 11408 3968
rect 11442 3792 11454 3968
rect 11396 3780 11454 3792
rect 11138 3550 11196 3562
rect 11138 3374 11150 3550
rect 11184 3374 11196 3550
rect 11138 3362 11196 3374
rect 11396 3550 11454 3562
rect 11396 3374 11408 3550
rect 11442 3374 11454 3550
rect 11396 3362 11454 3374
rect 11138 3132 11196 3144
rect 11138 2956 11150 3132
rect 11184 2956 11196 3132
rect 11138 2944 11196 2956
rect 11396 3132 11454 3144
rect 11396 2956 11408 3132
rect 11442 2956 11454 3132
rect 11396 2944 11454 2956
rect 11138 2714 11196 2726
rect 11138 2538 11150 2714
rect 11184 2538 11196 2714
rect 11138 2526 11196 2538
rect 11396 2714 11454 2726
rect 11396 2538 11408 2714
rect 11442 2538 11454 2714
rect 11396 2526 11454 2538
rect 11138 2296 11196 2308
rect 11138 2120 11150 2296
rect 11184 2120 11196 2296
rect 11138 2108 11196 2120
rect 11396 2296 11454 2308
rect 11396 2120 11408 2296
rect 11442 2120 11454 2296
rect 11396 2108 11454 2120
rect 11138 1878 11196 1890
rect 11138 1702 11150 1878
rect 11184 1702 11196 1878
rect 11138 1690 11196 1702
rect 11396 1878 11454 1890
rect 11396 1702 11408 1878
rect 11442 1702 11454 1878
rect 11396 1690 11454 1702
<< pdiff >>
rect 3338 4507 3396 4519
rect 3338 4131 3350 4507
rect 3384 4131 3396 4507
rect 3338 4119 3396 4131
rect 3596 4507 3654 4519
rect 3596 4131 3608 4507
rect 3642 4131 3654 4507
rect 3596 4119 3654 4131
rect 8158 4507 8216 4519
rect 8158 4131 8170 4507
rect 8204 4131 8216 4507
rect 8158 4119 8216 4131
rect 8416 4507 8474 4519
rect 8416 4131 8428 4507
rect 8462 4131 8474 4507
rect 8416 4119 8474 4131
rect 2638 3387 2696 3399
rect 2638 3011 2650 3387
rect 2684 3011 2696 3387
rect 2638 2999 2696 3011
rect 2896 3387 2954 3399
rect 2896 3011 2908 3387
rect 2942 3011 2954 3387
rect 2896 2999 2954 3011
rect 3158 2267 3216 2279
rect 3158 1891 3170 2267
rect 3204 1891 3216 2267
rect 3158 1879 3216 1891
rect 3416 2267 3474 2279
rect 3416 1891 3428 2267
rect 3462 1891 3474 2267
rect 3416 1879 3474 1891
rect 6538 2267 6596 2279
rect 6538 1891 6550 2267
rect 6584 1891 6596 2267
rect 6538 1879 6596 1891
rect 6796 2267 6854 2279
rect 6796 1891 6808 2267
rect 6842 1891 6854 2267
rect 6796 1879 6854 1891
<< ndiffc >>
rect 11150 4628 11184 4804
rect 11408 4628 11442 4804
rect 11150 4210 11184 4386
rect 11408 4210 11442 4386
rect 11150 3792 11184 3968
rect 11408 3792 11442 3968
rect 11150 3374 11184 3550
rect 11408 3374 11442 3550
rect 11150 2956 11184 3132
rect 11408 2956 11442 3132
rect 11150 2538 11184 2714
rect 11408 2538 11442 2714
rect 11150 2120 11184 2296
rect 11408 2120 11442 2296
rect 11150 1702 11184 1878
rect 11408 1702 11442 1878
<< pdiffc >>
rect 3350 4131 3384 4507
rect 3608 4131 3642 4507
rect 8170 4131 8204 4507
rect 8428 4131 8462 4507
rect 2650 3011 2684 3387
rect 2908 3011 2942 3387
rect 3170 1891 3204 2267
rect 3428 1891 3462 2267
rect 6550 1891 6584 2267
rect 6808 1891 6842 2267
<< psubdiff >>
rect 10686 5090 10710 5170
rect 10850 5090 10874 5170
rect 11036 4956 11132 4990
rect 11460 4956 11556 4990
rect 11036 4894 11070 4956
rect 11522 4894 11556 4956
rect 11036 1550 11070 1612
rect 11522 1550 11556 1612
rect 11036 1516 11132 1550
rect 11460 1516 11556 1550
<< nsubdiff >>
rect 3236 4668 3332 4702
rect 3660 4668 3756 4702
rect 3236 4606 3270 4668
rect 3722 4606 3756 4668
rect 3236 3970 3270 4032
rect 3722 3970 3756 4032
rect 3236 3936 3332 3970
rect 3660 3936 3756 3970
rect 8056 4668 8152 4702
rect 8480 4668 8576 4702
rect 8056 4606 8090 4668
rect 8542 4606 8576 4668
rect 8056 3970 8090 4032
rect 8542 3970 8576 4032
rect 8056 3936 8152 3970
rect 8480 3936 8576 3970
rect 2536 3548 2632 3582
rect 2960 3548 3056 3582
rect 2536 3486 2570 3548
rect 3022 3486 3056 3548
rect 2536 2850 2570 2912
rect 3022 2850 3056 2912
rect 2536 2816 2632 2850
rect 2960 2816 3056 2850
rect 3056 2428 3152 2462
rect 3480 2428 3576 2462
rect 3056 2366 3090 2428
rect 3542 2366 3576 2428
rect 3056 1730 3090 1792
rect 3542 1730 3576 1792
rect 3056 1696 3152 1730
rect 3480 1696 3576 1730
rect 6436 2428 6532 2462
rect 6860 2428 6956 2462
rect 6436 2366 6470 2428
rect 6922 2366 6956 2428
rect 6436 1730 6470 1792
rect 6922 1730 6956 1792
rect 6436 1696 6532 1730
rect 6860 1696 6956 1730
<< psubdiffcont >>
rect 10710 5090 10850 5170
rect 11132 4956 11460 4990
rect 11036 1612 11070 4894
rect 11522 1612 11556 4894
rect 11132 1516 11460 1550
<< nsubdiffcont >>
rect 3332 4668 3660 4702
rect 3236 4032 3270 4606
rect 3722 4032 3756 4606
rect 3332 3936 3660 3970
rect 8152 4668 8480 4702
rect 8056 4032 8090 4606
rect 8542 4032 8576 4606
rect 8152 3936 8480 3970
rect 2632 3548 2960 3582
rect 2536 2912 2570 3486
rect 3022 2912 3056 3486
rect 2632 2816 2960 2850
rect 3152 2428 3480 2462
rect 3056 1792 3090 2366
rect 3542 1792 3576 2366
rect 3152 1696 3480 1730
rect 6532 2428 6860 2462
rect 6436 1792 6470 2366
rect 6922 1792 6956 2366
rect 6532 1696 6860 1730
<< poly >>
rect 3396 4600 3596 4616
rect 3396 4566 3412 4600
rect 3580 4566 3596 4600
rect 3396 4519 3596 4566
rect 3396 4072 3596 4119
rect 3396 4038 3412 4072
rect 3580 4038 3596 4072
rect 3396 4022 3596 4038
rect 8216 4600 8416 4616
rect 8216 4566 8232 4600
rect 8400 4566 8416 4600
rect 8216 4519 8416 4566
rect 8216 4072 8416 4119
rect 8216 4038 8232 4072
rect 8400 4038 8416 4072
rect 8216 4022 8416 4038
rect 2696 3480 2896 3496
rect 2696 3446 2712 3480
rect 2880 3446 2896 3480
rect 2696 3399 2896 3446
rect 2696 2952 2896 2999
rect 2696 2918 2712 2952
rect 2880 2918 2896 2952
rect 2696 2902 2896 2918
rect 3216 2360 3416 2376
rect 3216 2326 3232 2360
rect 3400 2326 3416 2360
rect 3216 2279 3416 2326
rect 3216 1832 3416 1879
rect 3216 1798 3232 1832
rect 3400 1798 3416 1832
rect 3216 1782 3416 1798
rect 6596 2360 6796 2376
rect 6596 2326 6612 2360
rect 6780 2326 6796 2360
rect 6596 2279 6796 2326
rect 6596 1832 6796 1879
rect 6596 1798 6612 1832
rect 6780 1798 6796 1832
rect 6596 1782 6796 1798
rect 11196 4888 11396 4904
rect 11196 4854 11212 4888
rect 11380 4854 11396 4888
rect 11196 4816 11396 4854
rect 11196 4578 11396 4616
rect 11196 4544 11212 4578
rect 11380 4544 11396 4578
rect 11196 4528 11396 4544
rect 11196 4470 11396 4486
rect 11196 4436 11212 4470
rect 11380 4436 11396 4470
rect 11196 4398 11396 4436
rect 11196 4160 11396 4198
rect 11196 4126 11212 4160
rect 11380 4126 11396 4160
rect 11196 4110 11396 4126
rect 11196 4052 11396 4068
rect 11196 4018 11212 4052
rect 11380 4018 11396 4052
rect 11196 3980 11396 4018
rect 11196 3742 11396 3780
rect 11196 3708 11212 3742
rect 11380 3708 11396 3742
rect 11196 3692 11396 3708
rect 11196 3634 11396 3650
rect 11196 3600 11212 3634
rect 11380 3600 11396 3634
rect 11196 3562 11396 3600
rect 11196 3324 11396 3362
rect 11196 3290 11212 3324
rect 11380 3290 11396 3324
rect 11196 3274 11396 3290
rect 11196 3216 11396 3232
rect 11196 3182 11212 3216
rect 11380 3182 11396 3216
rect 11196 3144 11396 3182
rect 11196 2906 11396 2944
rect 11196 2872 11212 2906
rect 11380 2872 11396 2906
rect 11196 2856 11396 2872
rect 11196 2798 11396 2814
rect 11196 2764 11212 2798
rect 11380 2764 11396 2798
rect 11196 2726 11396 2764
rect 11196 2488 11396 2526
rect 11196 2454 11212 2488
rect 11380 2454 11396 2488
rect 11196 2438 11396 2454
rect 11196 2380 11396 2396
rect 11196 2346 11212 2380
rect 11380 2346 11396 2380
rect 11196 2308 11396 2346
rect 11196 2070 11396 2108
rect 11196 2036 11212 2070
rect 11380 2036 11396 2070
rect 11196 2020 11396 2036
rect 11196 1962 11396 1978
rect 11196 1928 11212 1962
rect 11380 1928 11396 1962
rect 11196 1890 11396 1928
rect 11196 1652 11396 1690
rect 11196 1618 11212 1652
rect 11380 1618 11396 1652
rect 11196 1602 11396 1618
<< polycont >>
rect 3412 4566 3580 4600
rect 3412 4038 3580 4072
rect 8232 4566 8400 4600
rect 8232 4038 8400 4072
rect 2712 3446 2880 3480
rect 2712 2918 2880 2952
rect 3232 2326 3400 2360
rect 3232 1798 3400 1832
rect 6612 2326 6780 2360
rect 6612 1798 6780 1832
rect 11212 4854 11380 4888
rect 11212 4544 11380 4578
rect 11212 4436 11380 4470
rect 11212 4126 11380 4160
rect 11212 4018 11380 4052
rect 11212 3708 11380 3742
rect 11212 3600 11380 3634
rect 11212 3290 11380 3324
rect 11212 3182 11380 3216
rect 11212 2872 11380 2906
rect 11212 2764 11380 2798
rect 11212 2454 11380 2488
rect 11212 2346 11380 2380
rect 11212 2036 11380 2070
rect 11212 1928 11380 1962
rect 11212 1618 11380 1652
<< locali >>
rect 11036 4894 11070 4990
rect 3236 4668 3332 4702
rect 3660 4668 3756 4702
rect 3236 4606 3270 4668
rect 3722 4606 3756 4668
rect 3396 4566 3412 4600
rect 3580 4566 3596 4600
rect 3350 4507 3384 4523
rect 3350 4115 3384 4131
rect 3608 4507 3642 4523
rect 3608 4115 3642 4131
rect 3396 4038 3412 4072
rect 3580 4038 3596 4072
rect 3236 3970 3270 4032
rect 3722 3970 3756 4032
rect 3236 3936 3332 3970
rect 3660 3936 3756 3970
rect 8056 4668 8152 4702
rect 8480 4668 8576 4702
rect 8056 4606 8090 4668
rect 8542 4606 8576 4668
rect 8216 4566 8232 4600
rect 8400 4566 8416 4600
rect 8170 4507 8204 4523
rect 8170 4115 8204 4131
rect 8428 4507 8462 4523
rect 8428 4115 8462 4131
rect 8216 4038 8232 4072
rect 8400 4038 8416 4072
rect 8056 3970 8090 4032
rect 8542 3970 8576 4032
rect 8056 3936 8152 3970
rect 8480 3936 8576 3970
rect 2536 3548 2632 3582
rect 2960 3548 3056 3582
rect 2536 3486 2570 3548
rect 3022 3486 3056 3548
rect 2696 3446 2712 3480
rect 2880 3446 2896 3480
rect 2650 3387 2684 3403
rect 2650 2995 2684 3011
rect 2908 3387 2942 3403
rect 2908 2995 2942 3011
rect 2696 2918 2712 2952
rect 2880 2918 2896 2952
rect 2536 2850 2570 2912
rect 3022 2850 3056 2912
rect 2536 2816 2632 2850
rect 2960 2816 3056 2850
rect 3056 2428 3152 2462
rect 3480 2428 3576 2462
rect 3056 2366 3090 2428
rect 3542 2366 3576 2428
rect 3216 2326 3232 2360
rect 3400 2326 3416 2360
rect 3170 2267 3204 2283
rect 3170 1875 3204 1891
rect 3428 2267 3462 2283
rect 3428 1875 3462 1891
rect 3216 1798 3232 1832
rect 3400 1798 3416 1832
rect 3056 1730 3090 1792
rect 3542 1730 3576 1792
rect 3056 1696 3152 1730
rect 3480 1696 3576 1730
rect 6436 2428 6532 2462
rect 6860 2428 6956 2462
rect 6436 2366 6470 2428
rect 6922 2366 6956 2428
rect 6596 2326 6612 2360
rect 6780 2326 6796 2360
rect 6550 2267 6584 2283
rect 6550 1875 6584 1891
rect 6808 2267 6842 2283
rect 6808 1875 6842 1891
rect 6596 1798 6612 1832
rect 6780 1798 6796 1832
rect 6436 1730 6470 1792
rect 6922 1730 6956 1792
rect 6436 1696 6532 1730
rect 6860 1696 6956 1730
rect 11522 4894 11556 4990
rect 11196 4854 11212 4888
rect 11380 4854 11396 4888
rect 11150 4804 11184 4820
rect 11150 4612 11184 4628
rect 11408 4804 11442 4820
rect 11408 4612 11442 4628
rect 11196 4544 11212 4578
rect 11380 4544 11396 4578
rect 11196 4436 11212 4470
rect 11380 4436 11396 4470
rect 11150 4386 11184 4402
rect 11150 4194 11184 4210
rect 11408 4386 11442 4402
rect 11408 4194 11442 4210
rect 11196 4126 11212 4160
rect 11380 4126 11396 4160
rect 11196 4018 11212 4052
rect 11380 4018 11396 4052
rect 11150 3968 11184 3984
rect 11150 3776 11184 3792
rect 11408 3968 11442 3984
rect 11408 3776 11442 3792
rect 11196 3708 11212 3742
rect 11380 3708 11396 3742
rect 11196 3600 11212 3634
rect 11380 3600 11396 3634
rect 11150 3550 11184 3566
rect 11150 3358 11184 3374
rect 11408 3550 11442 3566
rect 11408 3358 11442 3374
rect 11196 3290 11212 3324
rect 11380 3290 11396 3324
rect 11196 3182 11212 3216
rect 11380 3182 11396 3216
rect 11150 3132 11184 3148
rect 11150 2940 11184 2956
rect 11408 3132 11442 3148
rect 11408 2940 11442 2956
rect 11196 2872 11212 2906
rect 11380 2872 11396 2906
rect 11196 2764 11212 2798
rect 11380 2764 11396 2798
rect 11150 2714 11184 2730
rect 11150 2522 11184 2538
rect 11408 2714 11442 2730
rect 11408 2522 11442 2538
rect 11196 2454 11212 2488
rect 11380 2454 11396 2488
rect 11196 2346 11212 2380
rect 11380 2346 11396 2380
rect 11150 2296 11184 2312
rect 11150 2104 11184 2120
rect 11408 2296 11442 2312
rect 11408 2104 11442 2120
rect 11196 2036 11212 2070
rect 11380 2036 11396 2070
rect 11196 1928 11212 1962
rect 11380 1928 11396 1962
rect 11150 1878 11184 1894
rect 11150 1686 11184 1702
rect 11408 1878 11442 1894
rect 11408 1686 11442 1702
rect 11196 1618 11212 1652
rect 11380 1618 11396 1652
rect 11036 1550 11070 1612
rect 11522 1550 11556 1612
rect 11036 1516 11132 1550
rect 11460 1516 11556 1550
<< viali >>
rect 10690 5090 10710 5170
rect 10710 5090 10850 5170
rect 10850 5090 10870 5170
rect 11070 4956 11132 4990
rect 11132 4956 11460 4990
rect 11460 4956 11522 4990
rect 11212 4854 11380 4888
rect 11150 4628 11184 4804
rect 11408 4628 11442 4804
rect 11212 4544 11380 4578
rect 11212 4436 11380 4470
rect 11150 4210 11184 4386
rect 11408 4210 11442 4386
rect 11212 4126 11380 4160
rect 11212 4018 11380 4052
rect 11150 3792 11184 3968
rect 11408 3792 11442 3968
rect 11212 3708 11380 3742
rect 11212 3600 11380 3634
rect 11150 3374 11184 3550
rect 11408 3374 11442 3550
rect 11212 3290 11380 3324
rect 11212 3182 11380 3216
rect 11150 2956 11184 3132
rect 11408 2956 11442 3132
rect 11212 2872 11380 2906
rect 11212 2764 11380 2798
rect 11150 2538 11184 2714
rect 11408 2538 11442 2714
rect 11212 2454 11380 2488
rect 11212 2346 11380 2380
rect 11150 2120 11184 2296
rect 11408 2120 11442 2296
rect 11212 2036 11380 2070
rect 11212 1928 11380 1962
rect 11150 1702 11184 1878
rect 11408 1702 11442 1878
rect 11212 1618 11380 1652
<< metal1 >>
rect 4620 4960 4820 5340
rect 9960 5140 10160 5340
rect 9980 5080 10160 5140
rect 10660 5170 10880 5200
rect 10660 5090 10690 5170
rect 10870 5090 10880 5170
rect 10660 5080 10880 5090
rect 9160 5060 10880 5080
rect 9160 4980 9180 5060
rect 9260 4980 9320 5060
rect 9400 4980 9480 5060
rect 9560 4980 9660 5060
rect 9740 4980 9840 5060
rect 9920 4980 10020 5060
rect 10100 4980 10200 5060
rect 10280 4980 10380 5060
rect 10460 4980 10540 5060
rect 10620 4980 10720 5060
rect 10800 4980 10880 5060
rect 9160 4960 10880 4980
rect 11058 4990 11534 4996
rect 3080 4740 6200 4960
rect 11058 4956 11070 4990
rect 11522 4956 11534 4990
rect 11058 4950 11534 4956
rect 11200 4888 11392 4894
rect 11200 4854 11212 4888
rect 11380 4854 11392 4888
rect 11200 4848 11392 4854
rect 3080 2260 3360 4740
rect 4100 4440 4220 4740
rect 5600 4520 5720 4700
rect 5040 4500 5920 4520
rect 5040 4440 5840 4500
rect 5900 4440 5920 4500
rect 5820 4420 5920 4440
rect 6060 4400 6200 4740
rect 6700 4500 6900 4520
rect 7000 4500 7060 4700
rect 6700 4440 6720 4500
rect 6780 4440 6820 4500
rect 6880 4440 7600 4500
rect 6700 4420 6900 4440
rect 4480 4060 4640 4400
rect 5820 4300 5920 4320
rect 5320 4240 5840 4300
rect 5340 4180 5840 4240
rect 5900 4180 5920 4300
rect 5340 4160 5920 4180
rect 6460 4060 6620 4380
rect 6700 4300 6900 4320
rect 6700 4180 6720 4300
rect 6780 4180 6820 4300
rect 6880 4180 7340 4300
rect 6700 4160 7340 4180
rect 4260 4020 7560 4060
rect 4260 3840 9080 4020
rect 4100 3620 8820 3760
rect 4100 3380 4280 3620
rect 5740 3400 5800 3580
rect 5940 3400 6140 3420
rect 3520 3320 4280 3380
rect 4640 3340 5960 3400
rect 6020 3340 6060 3400
rect 6120 3340 6140 3400
rect 6240 3400 6300 3620
rect 7000 3400 7280 3420
rect 7340 3400 7400 3580
rect 6240 3340 6840 3400
rect 7000 3340 7020 3400
rect 7080 3340 7100 3400
rect 7160 3340 7200 3400
rect 7260 3340 8480 3400
rect 8660 3340 8820 3620
rect 4640 3320 6140 3340
rect 7000 3320 7280 3340
rect 7400 3320 8460 3340
rect 8660 3280 8680 3340
rect 8800 3280 8820 3340
rect 8660 3260 8820 3280
rect 8940 3340 9080 3840
rect 9160 3340 9260 4820
rect 9500 4720 9580 4800
rect 9500 4620 9580 4640
rect 9840 4720 9900 4820
rect 10140 4740 10220 4810
rect 9840 4640 9940 4720
rect 10140 4640 10220 4660
rect 9840 4590 10060 4640
rect 9310 4580 9480 4590
rect 9310 4520 9320 4580
rect 9470 4520 9480 4580
rect 9310 4510 9480 4520
rect 9840 4580 10120 4590
rect 9840 4520 9960 4580
rect 10110 4520 10120 4580
rect 9500 4300 9580 4380
rect 9500 4200 9580 4220
rect 9840 4300 9900 4520
rect 9950 4510 10120 4520
rect 10140 4360 10240 4380
rect 9840 4220 9940 4300
rect 10140 4220 10160 4360
rect 10220 4220 10240 4360
rect 9840 4170 10060 4220
rect 10140 4200 10240 4220
rect 9300 4160 9480 4170
rect 9300 4100 9310 4160
rect 9470 4100 9480 4160
rect 9300 4090 9480 4100
rect 9840 4160 10130 4170
rect 9840 4100 9970 4160
rect 10120 4100 10130 4160
rect 9500 3880 9580 3960
rect 9500 3780 9580 3800
rect 9840 3880 9900 4100
rect 9960 4090 10130 4100
rect 10140 3900 10220 3980
rect 9840 3800 9940 3880
rect 10140 3800 10220 3820
rect 9840 3750 10060 3800
rect 9300 3740 9480 3750
rect 9300 3680 9310 3740
rect 9470 3680 9480 3740
rect 9300 3670 9480 3680
rect 9840 3740 10120 3750
rect 9840 3680 9960 3740
rect 10110 3680 10120 3740
rect 9500 3480 9580 3560
rect 9500 3380 9580 3400
rect 9840 3480 9900 3680
rect 9950 3670 10120 3680
rect 10140 3480 10220 3560
rect 9840 3380 9940 3480
rect 10140 3380 10220 3400
rect 8940 3180 9260 3340
rect 9840 3330 10060 3380
rect 9300 3320 9480 3330
rect 9300 3260 9310 3320
rect 9470 3260 9480 3320
rect 9300 3250 9480 3260
rect 9840 3320 10120 3330
rect 9840 3260 9960 3320
rect 10110 3260 10120 3320
rect 4700 3160 4800 3180
rect 3760 3040 4720 3160
rect 4780 3040 4800 3160
rect 3760 3020 4800 3040
rect 4900 2960 5460 3180
rect 5940 3160 6140 3180
rect 5940 3040 5960 3160
rect 6020 3040 6060 3160
rect 6120 3040 6600 3160
rect 5940 3020 6600 3040
rect 7660 2960 8220 3180
rect 3540 2820 8420 2960
rect 5660 2520 5900 2820
rect 5660 2500 6380 2520
rect 4080 2320 6380 2500
rect 4280 2260 4640 2280
rect 3080 1880 4060 2260
rect 4280 2200 4500 2260
rect 4620 2200 4640 2260
rect 4280 2160 4640 2200
rect 5900 2260 6040 2280
rect 5900 2200 5960 2260
rect 6020 2200 6040 2260
rect 5900 2180 6040 2200
rect 4280 2100 4500 2160
rect 4620 2100 4640 2160
rect 4280 2060 4640 2100
rect 4280 2000 4500 2060
rect 4620 2000 4640 2060
rect 4280 1960 4640 2000
rect 4280 1900 4500 1960
rect 4620 1900 4640 1960
rect 5940 2160 6040 2180
rect 5940 2100 5960 2160
rect 6020 2100 6040 2160
rect 5940 2080 6040 2100
rect 5940 2020 5960 2080
rect 6020 2020 6040 2080
rect 5940 1980 6040 2020
rect 4280 1880 4640 1900
rect 3080 1660 3960 1880
rect 4740 1720 4900 1940
rect 5940 1920 5960 1980
rect 6020 1920 6040 1980
rect 5940 1900 6040 1920
rect 6120 2200 6380 2320
rect 6120 1900 9100 2200
rect 4740 1660 6060 1720
rect 3080 1500 6060 1660
rect 6120 1480 6380 1900
rect 7400 1560 7640 1580
rect 7400 1500 7420 1560
rect 7520 1500 7560 1560
rect 7620 1500 7640 1560
rect 7400 1480 7640 1500
rect 8860 1480 9100 1900
rect 9160 1680 9260 3180
rect 9500 3060 9580 3140
rect 9500 2960 9580 2980
rect 9840 3040 9900 3260
rect 9950 3250 10120 3260
rect 10140 3060 10220 3140
rect 9840 2960 9940 3040
rect 10140 2960 10220 2980
rect 9840 2920 10060 2960
rect 9310 2910 9480 2920
rect 9310 2850 9320 2910
rect 9470 2850 9480 2910
rect 9310 2840 9480 2850
rect 9840 2910 10120 2920
rect 9840 2850 9960 2910
rect 10110 2850 10120 2910
rect 9840 2840 10120 2850
rect 9500 2640 9580 2720
rect 9500 2540 9580 2560
rect 9840 2620 9900 2840
rect 10140 2640 10220 2720
rect 9840 2540 9940 2620
rect 10140 2540 10220 2560
rect 9840 2500 10060 2540
rect 9310 2490 9480 2500
rect 9310 2430 9320 2490
rect 9470 2430 9480 2490
rect 9310 2420 9480 2430
rect 9840 2490 10130 2500
rect 9840 2430 9970 2490
rect 10120 2430 10130 2490
rect 9840 2420 10130 2430
rect 9500 2220 9580 2300
rect 9500 2120 9580 2140
rect 9840 2200 9900 2420
rect 10140 2220 10220 2300
rect 9840 2120 9940 2200
rect 10140 2120 10220 2140
rect 9840 2080 10060 2120
rect 9310 2070 9480 2080
rect 9310 2010 9320 2070
rect 9470 2010 9480 2070
rect 9310 2000 9480 2010
rect 9840 2070 10130 2080
rect 9840 2010 9970 2070
rect 10120 2010 10130 2070
rect 9840 2000 10130 2010
rect 9500 1800 9580 1880
rect 9500 1700 9580 1720
rect 9840 1800 9900 2000
rect 10140 1800 10220 1880
rect 9840 1700 9940 1800
rect 10140 1700 10220 1720
rect 9840 1660 10060 1700
rect 9320 1650 9490 1660
rect 9320 1590 9330 1650
rect 9480 1590 9490 1650
rect 9320 1580 9490 1590
rect 9840 1650 10130 1660
rect 9840 1590 9970 1650
rect 10120 1590 10130 1650
rect 9840 1580 10130 1590
rect 10360 1480 10540 4820
rect 10780 4740 10860 4810
rect 10780 4640 10860 4660
rect 11144 4804 11190 4816
rect 11144 4628 11150 4804
rect 11184 4628 11190 4804
rect 11144 4616 11190 4628
rect 11402 4804 11448 4816
rect 11402 4628 11408 4804
rect 11442 4628 11448 4804
rect 11402 4616 11448 4628
rect 10590 4580 10760 4590
rect 10590 4520 10600 4580
rect 10750 4520 10760 4580
rect 11200 4578 11392 4584
rect 11200 4544 11212 4578
rect 11380 4544 11392 4578
rect 11200 4538 11392 4544
rect 10590 4510 10760 4520
rect 11200 4470 11392 4476
rect 11200 4436 11212 4470
rect 11380 4436 11392 4470
rect 11200 4430 11392 4436
rect 10780 4320 10860 4390
rect 10780 4220 10860 4240
rect 11144 4386 11190 4398
rect 11144 4210 11150 4386
rect 11184 4210 11190 4386
rect 11144 4198 11190 4210
rect 11402 4386 11448 4398
rect 11402 4210 11408 4386
rect 11442 4210 11448 4386
rect 11402 4198 11448 4210
rect 10590 4160 10760 4170
rect 10590 4100 10600 4160
rect 10750 4100 10760 4160
rect 11200 4160 11392 4166
rect 11200 4126 11212 4160
rect 11380 4126 11392 4160
rect 11200 4120 11392 4126
rect 10590 4090 10760 4100
rect 11200 4052 11392 4058
rect 11200 4018 11212 4052
rect 11380 4018 11392 4052
rect 11200 4012 11392 4018
rect 10780 3900 10860 3970
rect 10780 3800 10860 3820
rect 11144 3968 11190 3980
rect 11144 3792 11150 3968
rect 11184 3792 11190 3968
rect 11144 3780 11190 3792
rect 11402 3968 11448 3980
rect 11402 3792 11408 3968
rect 11442 3792 11448 3968
rect 11402 3780 11448 3792
rect 10590 3740 10760 3750
rect 10590 3680 10600 3740
rect 10750 3680 10760 3740
rect 11200 3742 11392 3748
rect 11200 3708 11212 3742
rect 11380 3708 11392 3742
rect 11200 3702 11392 3708
rect 10590 3670 10760 3680
rect 11200 3634 11392 3640
rect 11200 3600 11212 3634
rect 11380 3600 11392 3634
rect 11200 3594 11392 3600
rect 11144 3550 11190 3562
rect 10780 3480 10860 3550
rect 10780 3380 10860 3400
rect 11144 3374 11150 3550
rect 11184 3374 11190 3550
rect 11144 3362 11190 3374
rect 11402 3550 11448 3562
rect 11402 3374 11408 3550
rect 11442 3374 11448 3550
rect 11402 3362 11448 3374
rect 10590 3320 10760 3330
rect 10590 3260 10600 3320
rect 10750 3260 10760 3320
rect 11200 3324 11392 3330
rect 11200 3290 11212 3324
rect 11380 3290 11392 3324
rect 11200 3284 11392 3290
rect 10590 3250 10760 3260
rect 11200 3216 11392 3222
rect 11200 3182 11212 3216
rect 11380 3182 11392 3216
rect 11200 3176 11392 3182
rect 11144 3132 11190 3144
rect 10780 3060 10860 3130
rect 10780 2960 10860 2980
rect 11144 2956 11150 3132
rect 11184 2956 11190 3132
rect 11144 2944 11190 2956
rect 11402 3132 11448 3144
rect 11402 2956 11408 3132
rect 11442 2956 11448 3132
rect 11402 2944 11448 2956
rect 10590 2910 10760 2920
rect 10590 2850 10600 2910
rect 10750 2850 10760 2910
rect 11200 2906 11392 2912
rect 11200 2872 11212 2906
rect 11380 2872 11392 2906
rect 11200 2866 11392 2872
rect 10590 2840 10760 2850
rect 11200 2798 11392 2804
rect 11200 2764 11212 2798
rect 11380 2764 11392 2798
rect 11200 2758 11392 2764
rect 11144 2714 11190 2726
rect 10780 2640 10860 2710
rect 10780 2540 10860 2560
rect 11144 2538 11150 2714
rect 11184 2538 11190 2714
rect 11144 2526 11190 2538
rect 11402 2714 11448 2726
rect 11402 2538 11408 2714
rect 11442 2538 11448 2714
rect 11402 2526 11448 2538
rect 10590 2490 10760 2500
rect 10590 2430 10600 2490
rect 10750 2430 10760 2490
rect 11200 2488 11392 2494
rect 11200 2454 11212 2488
rect 11380 2454 11392 2488
rect 11200 2448 11392 2454
rect 10590 2420 10760 2430
rect 11200 2380 11392 2386
rect 11200 2346 11212 2380
rect 11380 2346 11392 2380
rect 11200 2340 11392 2346
rect 11144 2296 11190 2308
rect 10780 2220 10860 2290
rect 10780 2120 10860 2140
rect 11144 2120 11150 2296
rect 11184 2120 11190 2296
rect 11144 2108 11190 2120
rect 11402 2296 11448 2308
rect 11402 2120 11408 2296
rect 11442 2120 11448 2296
rect 11402 2108 11448 2120
rect 10600 2070 10770 2080
rect 10600 2010 10610 2070
rect 10760 2010 10770 2070
rect 11200 2070 11392 2076
rect 11200 2036 11212 2070
rect 11380 2036 11392 2070
rect 11200 2030 11392 2036
rect 10600 2000 10770 2010
rect 11200 1962 11392 1968
rect 11200 1928 11212 1962
rect 11380 1928 11392 1962
rect 11200 1922 11392 1928
rect 11144 1878 11190 1890
rect 10780 1800 10860 1870
rect 10780 1700 10860 1720
rect 11144 1702 11150 1878
rect 11184 1702 11190 1878
rect 11144 1690 11190 1702
rect 11402 1878 11448 1890
rect 11402 1702 11408 1878
rect 11442 1702 11448 1878
rect 11402 1690 11448 1702
rect 10590 1660 10760 1670
rect 10590 1600 10600 1660
rect 10750 1600 10760 1660
rect 11200 1652 11392 1658
rect 11200 1618 11212 1652
rect 11380 1618 11392 1652
rect 11200 1612 11392 1618
rect 10590 1590 10760 1600
rect 6140 1280 6340 1480
rect 7420 1280 7620 1480
rect 8860 1200 10540 1480
<< via1 >>
rect 9180 4980 9260 5060
rect 9320 4980 9400 5060
rect 9480 4980 9560 5060
rect 9660 4980 9740 5060
rect 9840 4980 9920 5060
rect 10020 4980 10100 5060
rect 10200 4980 10280 5060
rect 10380 4980 10460 5060
rect 10540 4980 10620 5060
rect 10720 4980 10800 5060
rect 5840 4440 5900 4500
rect 6720 4440 6780 4500
rect 6820 4440 6880 4500
rect 5840 4180 5900 4300
rect 6720 4180 6780 4300
rect 6820 4180 6880 4300
rect 5960 3340 6020 3400
rect 6060 3340 6120 3400
rect 7020 3340 7080 3400
rect 7100 3340 7160 3400
rect 7200 3340 7260 3400
rect 8680 3280 8800 3340
rect 9500 4640 9580 4720
rect 10140 4660 10220 4740
rect 9320 4520 9470 4580
rect 9960 4520 10110 4580
rect 9500 4220 9580 4300
rect 10160 4220 10220 4360
rect 9310 4100 9470 4160
rect 9970 4100 10120 4160
rect 9500 3800 9580 3880
rect 10140 3820 10220 3900
rect 9310 3680 9470 3740
rect 9960 3680 10110 3740
rect 9500 3400 9580 3480
rect 10140 3400 10220 3480
rect 9310 3260 9470 3320
rect 9960 3260 10110 3320
rect 4720 3040 4780 3160
rect 5960 3040 6020 3160
rect 6060 3040 6120 3160
rect 4500 2200 4620 2260
rect 5960 2200 6020 2260
rect 4500 2100 4620 2160
rect 4500 2000 4620 2060
rect 4500 1900 4620 1960
rect 5960 2100 6020 2160
rect 5960 2020 6020 2080
rect 5960 1920 6020 1980
rect 7420 1500 7520 1560
rect 7560 1500 7620 1560
rect 9500 2980 9580 3060
rect 10140 2980 10220 3060
rect 9320 2850 9470 2910
rect 9960 2850 10110 2910
rect 9500 2560 9580 2640
rect 10140 2560 10220 2640
rect 9320 2430 9470 2490
rect 9970 2430 10120 2490
rect 9500 2140 9580 2220
rect 10140 2140 10220 2220
rect 9320 2010 9470 2070
rect 9970 2010 10120 2070
rect 9500 1720 9580 1800
rect 10140 1720 10220 1800
rect 9330 1590 9480 1650
rect 9970 1590 10120 1650
rect 10780 4660 10860 4740
rect 10600 4520 10750 4580
rect 10780 4240 10860 4320
rect 10600 4100 10750 4160
rect 10780 3820 10860 3900
rect 10600 3680 10750 3740
rect 10780 3400 10860 3480
rect 10600 3260 10750 3320
rect 10780 2980 10860 3060
rect 10600 2850 10750 2910
rect 10780 2560 10860 2640
rect 10600 2430 10750 2490
rect 10780 2140 10860 2220
rect 10610 2010 10760 2070
rect 10780 1720 10860 1800
rect 10600 1600 10750 1660
<< metal2 >>
rect 9980 5080 10160 5140
rect 9160 5060 10880 5080
rect 9160 4980 9180 5060
rect 9260 4980 9320 5060
rect 9400 4980 9480 5060
rect 9560 4980 9660 5060
rect 9740 4980 9840 5060
rect 9920 4980 10020 5060
rect 10100 4980 10200 5060
rect 10280 4980 10380 5060
rect 10460 4980 10540 5060
rect 10620 4980 10720 5060
rect 10800 4980 10880 5060
rect 9160 4960 10880 4980
rect 10140 4810 10220 4819
rect 9500 4790 9580 4799
rect 4460 4580 6400 4680
rect 10140 4640 10220 4660
rect 10780 4810 10860 4819
rect 10780 4640 10860 4660
rect 9500 4620 9580 4640
rect 9310 4580 9480 4590
rect 9950 4580 10120 4590
rect 10590 4580 10760 4590
rect 4460 2260 4640 4580
rect 6260 4520 6400 4580
rect 9040 4520 9320 4580
rect 9470 4520 9960 4580
rect 10110 4520 10600 4580
rect 10750 4520 10760 4580
rect 5820 4500 6900 4520
rect 5820 4440 5840 4500
rect 5900 4440 6720 4500
rect 6780 4440 6820 4500
rect 6880 4440 6900 4500
rect 5820 4420 6900 4440
rect 5820 4300 5920 4320
rect 6700 4300 6900 4320
rect 5820 4180 5840 4300
rect 5900 4180 6720 4300
rect 6780 4180 6820 4300
rect 6880 4180 6900 4300
rect 5820 4160 6900 4180
rect 9040 4160 9100 4520
rect 9310 4510 9480 4520
rect 9950 4510 10120 4520
rect 10590 4510 10760 4520
rect 10780 4390 10860 4399
rect 9500 4370 9580 4379
rect 9500 4200 9580 4220
rect 10140 4360 10240 4380
rect 10140 4220 10160 4360
rect 10220 4220 10240 4360
rect 10780 4220 10860 4240
rect 10140 4200 10240 4220
rect 9300 4160 9480 4170
rect 9960 4160 10130 4170
rect 10590 4160 10760 4170
rect 6240 3820 6420 4160
rect 5100 3640 6420 3820
rect 9040 4100 9310 4160
rect 9470 4100 9970 4160
rect 10120 4100 10600 4160
rect 10750 4100 10980 4160
rect 9040 4080 10980 4100
rect 9040 3740 9100 4080
rect 10140 3970 10220 3979
rect 9500 3950 9580 3959
rect 10140 3800 10220 3820
rect 10780 3970 10860 3979
rect 10780 3800 10860 3820
rect 9500 3780 9580 3800
rect 9300 3740 9480 3750
rect 9950 3740 10120 3750
rect 10590 3740 10760 3750
rect 9040 3680 9310 3740
rect 9470 3680 9960 3740
rect 10110 3680 10600 3740
rect 10750 3680 10980 3740
rect 9040 3660 10980 3680
rect 4700 3160 4800 3180
rect 5100 3160 5320 3640
rect 5940 3400 6140 3420
rect 7000 3400 7280 3420
rect 5940 3340 5960 3400
rect 6020 3340 6060 3400
rect 6120 3340 7020 3400
rect 7080 3340 7100 3400
rect 7160 3340 7200 3400
rect 7260 3340 7440 3400
rect 5940 3320 7440 3340
rect 8660 3340 8820 3360
rect 9040 3340 9100 3660
rect 9500 3550 9580 3559
rect 9500 3380 9580 3400
rect 10140 3550 10220 3559
rect 10140 3380 10220 3400
rect 10780 3550 10860 3559
rect 10780 3380 10860 3400
rect 5940 3160 6140 3180
rect 4700 3040 4720 3160
rect 4780 3040 5960 3160
rect 6020 3040 6060 3160
rect 6120 3040 6140 3160
rect 4700 3020 6140 3040
rect 6480 2960 6680 3320
rect 8660 3280 8680 3340
rect 8800 3320 10760 3340
rect 8800 3280 9310 3320
rect 8660 3260 9310 3280
rect 9470 3260 9960 3320
rect 10110 3260 10600 3320
rect 10750 3260 10760 3320
rect 6220 2820 6680 2960
rect 9040 2920 9100 3260
rect 9300 3250 9480 3260
rect 9950 3250 10120 3260
rect 10590 3250 10760 3260
rect 9500 3130 9580 3139
rect 9500 2960 9580 2980
rect 10140 3130 10220 3139
rect 10140 2960 10220 2980
rect 10780 3130 10860 3139
rect 10780 2960 10860 2980
rect 9040 2910 10980 2920
rect 9040 2850 9320 2910
rect 9470 2850 9960 2910
rect 10110 2850 10600 2910
rect 10750 2850 10980 2910
rect 9040 2840 10980 2850
rect 6240 2280 6440 2820
rect 9040 2500 9100 2840
rect 9500 2710 9580 2719
rect 9500 2540 9580 2560
rect 10140 2710 10220 2719
rect 10140 2540 10220 2560
rect 10780 2710 10860 2719
rect 10780 2540 10860 2560
rect 9040 2490 10980 2500
rect 9040 2430 9320 2490
rect 9470 2430 9970 2490
rect 10120 2430 10600 2490
rect 10750 2430 10980 2490
rect 9040 2420 10980 2430
rect 4460 2200 4500 2260
rect 4620 2200 4640 2260
rect 4460 2160 4640 2200
rect 4460 2100 4500 2160
rect 4620 2100 4640 2160
rect 4460 2060 4640 2100
rect 4460 2000 4500 2060
rect 4620 2000 4640 2060
rect 4460 1960 4640 2000
rect 4460 1900 4500 1960
rect 4620 1900 4640 1960
rect 5940 2260 7640 2280
rect 5940 2200 5960 2260
rect 6020 2200 7640 2260
rect 5940 2160 7640 2200
rect 5940 2100 5960 2160
rect 6020 2100 7640 2160
rect 5940 2080 7640 2100
rect 5940 2020 5960 2080
rect 6020 2020 7640 2080
rect 5940 1980 7640 2020
rect 5940 1920 5960 1980
rect 6020 1920 7640 1980
rect 5940 1900 7640 1920
rect 4460 1880 4640 1900
rect 7400 1560 7640 1900
rect 9040 2080 9100 2420
rect 9500 2290 9580 2299
rect 9500 2120 9580 2140
rect 10140 2290 10220 2299
rect 10140 2120 10220 2140
rect 10780 2290 10860 2299
rect 10780 2120 10860 2140
rect 9040 2070 10980 2080
rect 9040 2010 9320 2070
rect 9470 2010 9970 2070
rect 10120 2010 10610 2070
rect 10760 2010 10980 2070
rect 9040 2000 10980 2010
rect 9040 1660 9100 2000
rect 9500 1870 9580 1879
rect 9500 1700 9580 1720
rect 10140 1870 10220 1879
rect 10140 1700 10220 1720
rect 10780 1870 10860 1879
rect 10780 1700 10860 1720
rect 10590 1660 10760 1670
rect 9040 1650 10600 1660
rect 9040 1590 9330 1650
rect 9480 1590 9970 1650
rect 10120 1600 10600 1650
rect 10750 1600 10980 1660
rect 10120 1590 10980 1600
rect 9040 1580 10980 1590
rect 7400 1500 7420 1560
rect 7520 1500 7560 1560
rect 7620 1500 7640 1560
rect 7400 1480 7640 1500
<< via2 >>
rect 9180 4980 9260 5060
rect 9320 4980 9400 5060
rect 9480 4980 9560 5060
rect 9660 4980 9740 5060
rect 9840 4980 9920 5060
rect 10020 4980 10100 5060
rect 10200 4980 10280 5060
rect 10380 4980 10460 5060
rect 10540 4980 10620 5060
rect 10720 4980 10800 5060
rect 9500 4720 9580 4790
rect 9500 4640 9580 4720
rect 10140 4740 10220 4810
rect 10140 4660 10220 4740
rect 10780 4740 10860 4810
rect 10780 4660 10860 4740
rect 9500 4300 9580 4370
rect 9500 4220 9580 4300
rect 10160 4220 10220 4360
rect 10780 4320 10860 4390
rect 10780 4240 10860 4320
rect 9500 3880 9580 3950
rect 9500 3800 9580 3880
rect 10140 3900 10220 3970
rect 10140 3820 10220 3900
rect 10780 3900 10860 3970
rect 10780 3820 10860 3900
rect 9500 3480 9580 3550
rect 9500 3400 9580 3480
rect 10140 3480 10220 3550
rect 10140 3400 10220 3480
rect 10780 3480 10860 3550
rect 10780 3400 10860 3480
rect 9500 3060 9580 3130
rect 9500 2980 9580 3060
rect 10140 3060 10220 3130
rect 10140 2980 10220 3060
rect 10780 3060 10860 3130
rect 10780 2980 10860 3060
rect 9500 2640 9580 2710
rect 9500 2560 9580 2640
rect 10140 2640 10220 2710
rect 10140 2560 10220 2640
rect 10780 2640 10860 2710
rect 10780 2560 10860 2640
rect 9500 2220 9580 2290
rect 9500 2140 9580 2220
rect 10140 2220 10220 2290
rect 10140 2140 10220 2220
rect 10780 2220 10860 2290
rect 10780 2140 10860 2220
rect 9500 1800 9580 1870
rect 9500 1720 9580 1800
rect 10140 1800 10220 1870
rect 10140 1720 10220 1800
rect 10780 1800 10860 1870
rect 10780 1720 10860 1800
<< metal3 >>
rect 9980 5080 10160 5140
rect 9160 5060 10880 5080
rect 9160 4980 9180 5060
rect 9260 4980 9320 5060
rect 9400 4980 9480 5060
rect 9560 4980 9660 5060
rect 9740 4980 9840 5060
rect 9920 4980 10020 5060
rect 10100 4980 10200 5060
rect 10280 4980 10380 5060
rect 10460 4980 10540 5060
rect 10620 4980 10720 5060
rect 10800 5000 10880 5060
rect 10800 4980 10920 5000
rect 9160 4960 10920 4980
rect 9520 4795 9660 4960
rect 10140 4815 10280 4960
rect 10780 4815 10920 4960
rect 9495 4790 9660 4795
rect 9495 4640 9500 4790
rect 9580 4640 9660 4790
rect 10135 4810 10280 4815
rect 10135 4660 10140 4810
rect 10220 4660 10280 4810
rect 10135 4655 10280 4660
rect 10775 4810 10920 4815
rect 10775 4660 10780 4810
rect 10860 4660 10920 4810
rect 10775 4655 10920 4660
rect 9495 4635 9660 4640
rect 9500 4620 9660 4635
rect 9520 4375 9660 4620
rect 9495 4370 9660 4375
rect 9495 4220 9500 4370
rect 9580 4220 9660 4370
rect 9495 4215 9660 4220
rect 9500 4200 9660 4215
rect 9520 3955 9660 4200
rect 10140 4360 10280 4655
rect 10780 4395 10920 4655
rect 10140 4220 10160 4360
rect 10220 4220 10280 4360
rect 10775 4390 10920 4395
rect 10775 4240 10780 4390
rect 10860 4240 10920 4390
rect 10775 4235 10920 4240
rect 10140 3975 10280 4220
rect 10780 3975 10920 4235
rect 9495 3950 9660 3955
rect 9495 3800 9500 3950
rect 9580 3800 9660 3950
rect 10135 3970 10280 3975
rect 10135 3820 10140 3970
rect 10220 3820 10280 3970
rect 10135 3815 10280 3820
rect 10775 3970 10920 3975
rect 10775 3820 10780 3970
rect 10860 3820 10920 3970
rect 10775 3815 10920 3820
rect 9495 3795 9660 3800
rect 9500 3780 9660 3795
rect 9520 3555 9660 3780
rect 10140 3555 10280 3815
rect 10780 3555 10920 3815
rect 9495 3550 9660 3555
rect 9495 3400 9500 3550
rect 9580 3400 9660 3550
rect 9495 3395 9660 3400
rect 10135 3550 10280 3555
rect 10135 3400 10140 3550
rect 10220 3400 10280 3550
rect 10135 3395 10280 3400
rect 10775 3550 10920 3555
rect 10775 3400 10780 3550
rect 10860 3400 10920 3550
rect 10775 3395 10920 3400
rect 9500 3380 9660 3395
rect 9520 3135 9660 3380
rect 10140 3135 10280 3395
rect 10780 3135 10920 3395
rect 9495 3130 9660 3135
rect 9495 2980 9500 3130
rect 9580 2980 9660 3130
rect 9495 2975 9660 2980
rect 10135 3130 10280 3135
rect 10135 2980 10140 3130
rect 10220 2980 10280 3130
rect 10135 2975 10280 2980
rect 10775 3130 10920 3135
rect 10775 2980 10780 3130
rect 10860 2980 10920 3130
rect 10775 2975 10920 2980
rect 9500 2960 9660 2975
rect 9520 2715 9660 2960
rect 10140 2715 10280 2975
rect 10780 2715 10920 2975
rect 9495 2710 9660 2715
rect 9495 2560 9500 2710
rect 9580 2560 9660 2710
rect 9495 2555 9660 2560
rect 10135 2710 10280 2715
rect 10135 2560 10140 2710
rect 10220 2560 10280 2710
rect 10135 2555 10280 2560
rect 10775 2710 10920 2715
rect 10775 2560 10780 2710
rect 10860 2560 10920 2710
rect 10775 2555 10920 2560
rect 9500 2540 9660 2555
rect 9520 2295 9660 2540
rect 10140 2295 10280 2555
rect 10780 2295 10920 2555
rect 9495 2290 9660 2295
rect 9495 2140 9500 2290
rect 9580 2140 9660 2290
rect 9495 2135 9660 2140
rect 10135 2290 10280 2295
rect 10135 2140 10140 2290
rect 10220 2140 10280 2290
rect 10135 2135 10280 2140
rect 10775 2290 10920 2295
rect 10775 2140 10780 2290
rect 10860 2140 10920 2290
rect 10775 2135 10920 2140
rect 9500 2120 9660 2135
rect 9520 1875 9660 2120
rect 10140 1875 10280 2135
rect 10780 1875 10920 2135
rect 9495 1870 9660 1875
rect 9495 1720 9500 1870
rect 9580 1720 9660 1870
rect 9495 1715 9660 1720
rect 10135 1870 10280 1875
rect 10135 1720 10140 1870
rect 10220 1720 10280 1870
rect 10135 1715 10280 1720
rect 10775 1870 10920 1875
rect 10775 1720 10780 1870
rect 10860 1720 10920 1870
rect 10775 1715 10920 1720
rect 9500 1700 9660 1715
rect 10140 1700 10280 1715
rect 10780 1700 10920 1715
use sky130_fd_pr__nfet_01v8_SXQYJB  XN3
timestamp 1657052488
transform 1 0 10676 0 1 3253
box -296 -1773 296 1773
use sky130_fd_pr__pfet_01v8_8CLM97  XP2
timestamp 1657122734
transform 1 0 7325 0 1 4319
box -425 -419 425 419
use sky130_fd_pr__pfet_01v8_82U688  XP4
timestamp 1657127204
transform 1 0 5436 0 1 2079
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_8CLZW6  XP6
timestamp 1657122734
transform 1 0 5183 0 1 3199
box -683 -419 683 419
use sky130_fd_pr__nfet_01v8_SXQYJB  sky130_fd_pr__nfet_01v8_SXQYJB_0
timestamp 1657052488
transform 1 0 10036 0 1 3253
box -296 -1773 296 1773
use sky130_fd_pr__nfet_01v8_SXQYJB  sky130_fd_pr__nfet_01v8_SXQYJB_1
timestamp 1657052488
transform 1 0 9396 0 1 3253
box -296 -1773 296 1773
use sky130_fd_pr__pfet_01v8_3P9HCE  sky130_fd_pr__pfet_01v8_3P9HCE_0
timestamp 1657122734
transform 1 0 6565 0 1 3199
box -425 -419 425 419
use sky130_fd_pr__pfet_01v8_8CLK97  sky130_fd_pr__pfet_01v8_8CLK97_0
timestamp 1657122734
transform 1 0 4356 0 1 4319
box -296 -419 296 419
use sky130_fd_pr__pfet_01v8_8CLK97  sky130_fd_pr__pfet_01v8_8CLK97_1
timestamp 1657122734
transform 1 0 6336 0 1 4319
box -296 -419 296 419
use sky130_fd_pr__pfet_01v8_8CLM97  sky130_fd_pr__pfet_01v8_8CLM97_0
timestamp 1657122734
transform 1 0 5345 0 1 4319
box -425 -419 425 419
use sky130_fd_pr__pfet_01v8_8CLZW6  sky130_fd_pr__pfet_01v8_8CLZW6_0
timestamp 1657122734
transform 1 0 7943 0 1 3199
box -683 -419 683 419
use sky130_fd_pr__pfet_01v8_37ZGCE  sky130_fd_pr__pfet_01v8_37ZGCE_0
timestamp 1657122734
transform 1 0 3785 0 1 3199
box -425 -419 425 419
use sky130_fd_pr__pfet_01v8_G8PMZT  sky130_fd_pr__pfet_01v8_G8PMZT_0
timestamp 1657052488
transform 1 0 4176 0 1 2079
box -296 -419 296 419
<< labels >>
flabel metal2 5820 3760 5820 3760 0 FreeSans 800 0 0 0 c
flabel metal1 8500 3640 8520 3660 0 FreeSans 800 0 0 0 b
flabel metal1 4620 5140 4820 5340 0 FreeSans 1600 0 0 0 vd
port 0 nsew
flabel metal1 9960 5140 10160 5340 0 FreeSans 1600 0 0 0 gnd
port 3 nsew
flabel metal2 4540 3760 4540 3760 0 FreeSans 800 0 0 0 d
flabel metal1 6980 3860 6980 3860 0 FreeSans 800 0 0 0 a
flabel metal1 7420 1280 7620 1480 0 FreeSans 1600 0 0 0 vts
port 1 nsew
flabel metal1 6140 1280 6340 1480 0 FreeSans 1600 0 0 0 vtd
port 2 nsew
<< end >>
