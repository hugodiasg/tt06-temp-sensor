magic
tech sky130A
magscale 1 2
timestamp 1708779589
<< metal2 >>
rect 9820 39240 10100 39250
rect 10100 38900 22540 39240
rect 9820 38880 22540 38900
rect 18050 34980 21760 35000
rect 18050 34800 18060 34980
rect 18260 34800 21760 34980
rect 18050 34780 21760 34800
rect 19280 34380 21720 34400
rect 19280 34220 19300 34380
rect 19460 34220 21720 34380
rect 19280 34200 21720 34220
rect 20640 26260 21680 26280
rect 20640 26100 20660 26260
rect 20820 26100 21680 26260
rect 20640 26080 21680 26100
rect 20640 25660 21780 25680
rect 20640 25500 20660 25660
rect 20820 25500 21780 25660
rect 20640 25480 21780 25500
rect 17600 25320 21600 25340
rect 17600 25160 17620 25320
rect 17780 25160 21600 25320
rect 17600 25140 21600 25160
rect 200 25080 480 25090
rect 190 24860 200 25080
rect 480 24860 21630 25080
rect 200 24850 480 24860
<< via2 >>
rect 9820 38900 10100 39240
rect 18060 34800 18260 34980
rect 19300 34220 19460 34380
rect 20660 26100 20820 26260
rect 20660 25500 20820 25660
rect 17620 25160 17780 25320
rect 200 24860 480 25080
<< metal3 >>
rect 17600 44620 17800 44660
rect 17600 44480 17620 44620
rect 17780 44480 17800 44620
rect 9810 39240 10110 39245
rect 9810 38900 9820 39240
rect 10100 38900 10110 39240
rect 9810 38895 10110 38900
rect 17600 25320 17800 44480
rect 20640 44500 20840 44520
rect 20640 44340 20660 44500
rect 20820 44340 20840 44500
rect 17600 25160 17620 25320
rect 17780 25160 17800 25320
rect 17600 25140 17800 25160
rect 18050 34980 18270 35000
rect 18050 34800 18060 34980
rect 18260 34800 18270 34980
rect 190 25080 490 25085
rect 190 24860 200 25080
rect 480 24860 490 25080
rect 190 24855 490 24860
rect 18050 1020 18270 34800
rect 18050 840 18060 1020
rect 18260 840 18270 1020
rect 18050 810 18270 840
rect 19280 34380 19480 34400
rect 19280 34220 19300 34380
rect 19460 34220 19480 34380
rect 19280 980 19480 34220
rect 20640 26260 20840 44340
rect 20640 26100 20660 26260
rect 20820 26100 20840 26260
rect 20640 26080 20840 26100
rect 20640 25660 20840 25680
rect 20640 25500 20660 25660
rect 20820 25500 20840 25660
rect 20640 3540 20840 25500
rect 20640 3380 20660 3540
rect 20820 3380 20840 3540
rect 20640 3360 20840 3380
rect 26860 3540 27060 3560
rect 26860 3380 26880 3540
rect 27040 3380 27060 3540
rect 19280 820 19300 980
rect 19460 820 19480 980
rect 26860 1100 27060 3380
rect 31000 1920 31440 32480
rect 31000 1560 31040 1920
rect 31400 1560 31440 1920
rect 31000 1520 31440 1560
rect 26860 940 26880 1100
rect 27040 940 27060 1100
rect 26860 920 27060 940
rect 19280 800 19480 820
<< via3 >>
rect 17620 44480 17780 44620
rect 9820 38900 10100 39240
rect 20660 44340 20820 44500
rect 200 24860 480 25080
rect 18060 840 18260 1020
rect 20660 3380 20820 3540
rect 26880 3380 27040 3540
rect 19300 820 19460 980
rect 31040 1560 31400 1920
rect 26880 940 27040 1100
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44820 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 17600 44620 17800 44820
rect 17600 44480 17620 44620
rect 17780 44480 17800 44620
rect 30974 44520 31034 45152
rect 31710 44952 31770 45152
rect 17600 44460 17800 44480
rect 20640 44500 31100 44520
rect 20640 44340 20660 44500
rect 20820 44340 31100 44500
rect 20640 44320 31100 44340
rect 200 25081 500 44152
rect 199 25080 500 25081
rect 199 24860 200 25080
rect 480 24860 500 25080
rect 199 24859 500 24860
rect 200 1000 500 24859
rect 9800 39241 10100 44152
rect 9800 39240 10101 39241
rect 9800 38900 9820 39240
rect 10100 38900 10101 39240
rect 9800 38899 10101 38900
rect 9800 1000 10100 38899
rect 20640 3540 27060 3560
rect 20640 3380 20660 3540
rect 20820 3380 26880 3540
rect 27040 3380 27060 3540
rect 20640 3360 27060 3380
rect 31000 1920 31440 1960
rect 31000 1560 31040 1920
rect 31400 1560 31440 1920
rect 26860 1100 27060 1120
rect 18050 1020 18270 1030
rect 18050 840 18060 1020
rect 18260 840 18270 1020
rect 18050 530 18270 840
rect 19280 980 22620 1000
rect 19280 820 19300 980
rect 19460 820 22620 980
rect 19280 800 22620 820
rect 26860 940 26880 1100
rect 27040 940 27060 1100
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 530
rect 22480 0 22600 800
rect 26860 500 27060 940
rect 31000 720 31440 1560
rect 26896 0 27016 500
rect 31312 0 31432 720
use device_without_rf  device_without_rf_0
timestamp 1708740906
transform 0 1 23870 -1 0 39352
box -62 -2580 29620 7540
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
