** sch_path: /home/hugodg/projects-sky130/temp-sensor/sensor/xschem/nmos_tb-dc.sch
**.subckt nmos_tb-dc
Va in GND 0.1
V2 out GND 1.8
XM1 GND in out out sky130_fd_pr__pfet_01v8 L=5 W=9.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.dc Va -2 2 0.001V
.control
run
set color0=white
set color1=black

let zout= out/(-i(v2))
let id=-I(v2)
plot zout
plot ph(zout)
plot id
*plot id xlimit 2.5 3.5 ylimit 0m 2m
.endc


.lib /home/hugodg/sky130_workspace/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
