magic
tech sky130A
magscale 1 2
timestamp 1656710231
<< pwell >>
rect -296 -1773 296 1773
<< nmos >>
rect -100 1363 100 1563
rect -100 945 100 1145
rect -100 527 100 727
rect -100 109 100 309
rect -100 -309 100 -109
rect -100 -727 100 -527
rect -100 -1145 100 -945
rect -100 -1563 100 -1363
<< ndiff >>
rect -158 1551 -100 1563
rect -158 1375 -146 1551
rect -112 1375 -100 1551
rect -158 1363 -100 1375
rect 100 1551 158 1563
rect 100 1375 112 1551
rect 146 1375 158 1551
rect 100 1363 158 1375
rect -158 1133 -100 1145
rect -158 957 -146 1133
rect -112 957 -100 1133
rect -158 945 -100 957
rect 100 1133 158 1145
rect 100 957 112 1133
rect 146 957 158 1133
rect 100 945 158 957
rect -158 715 -100 727
rect -158 539 -146 715
rect -112 539 -100 715
rect -158 527 -100 539
rect 100 715 158 727
rect 100 539 112 715
rect 146 539 158 715
rect 100 527 158 539
rect -158 297 -100 309
rect -158 121 -146 297
rect -112 121 -100 297
rect -158 109 -100 121
rect 100 297 158 309
rect 100 121 112 297
rect 146 121 158 297
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -297 -146 -121
rect -112 -297 -100 -121
rect -158 -309 -100 -297
rect 100 -121 158 -109
rect 100 -297 112 -121
rect 146 -297 158 -121
rect 100 -309 158 -297
rect -158 -539 -100 -527
rect -158 -715 -146 -539
rect -112 -715 -100 -539
rect -158 -727 -100 -715
rect 100 -539 158 -527
rect 100 -715 112 -539
rect 146 -715 158 -539
rect 100 -727 158 -715
rect -158 -957 -100 -945
rect -158 -1133 -146 -957
rect -112 -1133 -100 -957
rect -158 -1145 -100 -1133
rect 100 -957 158 -945
rect 100 -1133 112 -957
rect 146 -1133 158 -957
rect 100 -1145 158 -1133
rect -158 -1375 -100 -1363
rect -158 -1551 -146 -1375
rect -112 -1551 -100 -1375
rect -158 -1563 -100 -1551
rect 100 -1375 158 -1363
rect 100 -1551 112 -1375
rect 146 -1551 158 -1375
rect 100 -1563 158 -1551
<< ndiffc >>
rect -146 1375 -112 1551
rect 112 1375 146 1551
rect -146 957 -112 1133
rect 112 957 146 1133
rect -146 539 -112 715
rect 112 539 146 715
rect -146 121 -112 297
rect 112 121 146 297
rect -146 -297 -112 -121
rect 112 -297 146 -121
rect -146 -715 -112 -539
rect 112 -715 146 -539
rect -146 -1133 -112 -957
rect 112 -1133 146 -957
rect -146 -1551 -112 -1375
rect 112 -1551 146 -1375
<< psubdiff >>
rect -260 1703 -164 1737
rect 164 1703 260 1737
rect -260 1641 -226 1703
rect 226 1641 260 1703
rect -260 -1703 -226 -1641
rect 226 -1703 260 -1641
rect -260 -1737 -164 -1703
rect 164 -1737 260 -1703
<< psubdiffcont >>
rect -164 1703 164 1737
rect -260 -1641 -226 1641
rect 226 -1641 260 1641
rect -164 -1737 164 -1703
<< poly >>
rect -100 1635 100 1651
rect -100 1601 -84 1635
rect 84 1601 100 1635
rect -100 1563 100 1601
rect -100 1325 100 1363
rect -100 1291 -84 1325
rect 84 1291 100 1325
rect -100 1275 100 1291
rect -100 1217 100 1233
rect -100 1183 -84 1217
rect 84 1183 100 1217
rect -100 1145 100 1183
rect -100 907 100 945
rect -100 873 -84 907
rect 84 873 100 907
rect -100 857 100 873
rect -100 799 100 815
rect -100 765 -84 799
rect 84 765 100 799
rect -100 727 100 765
rect -100 489 100 527
rect -100 455 -84 489
rect 84 455 100 489
rect -100 439 100 455
rect -100 381 100 397
rect -100 347 -84 381
rect 84 347 100 381
rect -100 309 100 347
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -347 100 -309
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -397 100 -381
rect -100 -455 100 -439
rect -100 -489 -84 -455
rect 84 -489 100 -455
rect -100 -527 100 -489
rect -100 -765 100 -727
rect -100 -799 -84 -765
rect 84 -799 100 -765
rect -100 -815 100 -799
rect -100 -873 100 -857
rect -100 -907 -84 -873
rect 84 -907 100 -873
rect -100 -945 100 -907
rect -100 -1183 100 -1145
rect -100 -1217 -84 -1183
rect 84 -1217 100 -1183
rect -100 -1233 100 -1217
rect -100 -1291 100 -1275
rect -100 -1325 -84 -1291
rect 84 -1325 100 -1291
rect -100 -1363 100 -1325
rect -100 -1601 100 -1563
rect -100 -1635 -84 -1601
rect 84 -1635 100 -1601
rect -100 -1651 100 -1635
<< polycont >>
rect -84 1601 84 1635
rect -84 1291 84 1325
rect -84 1183 84 1217
rect -84 873 84 907
rect -84 765 84 799
rect -84 455 84 489
rect -84 347 84 381
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -381 84 -347
rect -84 -489 84 -455
rect -84 -799 84 -765
rect -84 -907 84 -873
rect -84 -1217 84 -1183
rect -84 -1325 84 -1291
rect -84 -1635 84 -1601
<< locali >>
rect -260 1703 -164 1737
rect 164 1703 260 1737
rect -260 1641 -226 1703
rect 226 1641 260 1703
rect -100 1601 -84 1635
rect 84 1601 100 1635
rect -146 1551 -112 1567
rect -146 1359 -112 1375
rect 112 1551 146 1567
rect 112 1359 146 1375
rect -100 1291 -84 1325
rect 84 1291 100 1325
rect -100 1183 -84 1217
rect 84 1183 100 1217
rect -146 1133 -112 1149
rect -146 941 -112 957
rect 112 1133 146 1149
rect 112 941 146 957
rect -100 873 -84 907
rect 84 873 100 907
rect -100 765 -84 799
rect 84 765 100 799
rect -146 715 -112 731
rect -146 523 -112 539
rect 112 715 146 731
rect 112 523 146 539
rect -100 455 -84 489
rect 84 455 100 489
rect -100 347 -84 381
rect 84 347 100 381
rect -146 297 -112 313
rect -146 105 -112 121
rect 112 297 146 313
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -313 -112 -297
rect 112 -121 146 -105
rect 112 -313 146 -297
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -489 -84 -455
rect 84 -489 100 -455
rect -146 -539 -112 -523
rect -146 -731 -112 -715
rect 112 -539 146 -523
rect 112 -731 146 -715
rect -100 -799 -84 -765
rect 84 -799 100 -765
rect -100 -907 -84 -873
rect 84 -907 100 -873
rect -146 -957 -112 -941
rect -146 -1149 -112 -1133
rect 112 -957 146 -941
rect 112 -1149 146 -1133
rect -100 -1217 -84 -1183
rect 84 -1217 100 -1183
rect -100 -1325 -84 -1291
rect 84 -1325 100 -1291
rect -146 -1375 -112 -1359
rect -146 -1567 -112 -1551
rect 112 -1375 146 -1359
rect 112 -1567 146 -1551
rect -100 -1635 -84 -1601
rect 84 -1635 100 -1601
rect -260 -1737 -226 -1641
rect 226 -1737 260 -1641
<< viali >>
rect -84 1601 84 1635
rect -146 1375 -112 1551
rect 112 1375 146 1551
rect -84 1291 84 1325
rect -84 1183 84 1217
rect -146 957 -112 1133
rect 112 957 146 1133
rect -84 873 84 907
rect -84 765 84 799
rect -146 539 -112 715
rect 112 539 146 715
rect -84 455 84 489
rect -84 347 84 381
rect -146 121 -112 297
rect 112 121 146 297
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -297 -112 -121
rect 112 -297 146 -121
rect -84 -381 84 -347
rect -84 -489 84 -455
rect -146 -715 -112 -539
rect 112 -715 146 -539
rect -84 -799 84 -765
rect -84 -907 84 -873
rect -146 -1133 -112 -957
rect 112 -1133 146 -957
rect -84 -1217 84 -1183
rect -84 -1325 84 -1291
rect -146 -1551 -112 -1375
rect 112 -1551 146 -1375
rect -84 -1635 84 -1601
rect -226 -1737 -164 -1703
rect -164 -1737 164 -1703
rect 164 -1737 226 -1703
<< metal1 >>
rect -96 1635 96 1641
rect -96 1601 -84 1635
rect 84 1601 96 1635
rect -96 1595 96 1601
rect -152 1551 -106 1563
rect -152 1375 -146 1551
rect -112 1375 -106 1551
rect -152 1363 -106 1375
rect 106 1551 152 1563
rect 106 1375 112 1551
rect 146 1375 152 1551
rect 106 1363 152 1375
rect -96 1325 96 1331
rect -96 1291 -84 1325
rect 84 1291 96 1325
rect -96 1285 96 1291
rect -96 1217 96 1223
rect -96 1183 -84 1217
rect 84 1183 96 1217
rect -96 1177 96 1183
rect -152 1133 -106 1145
rect -152 957 -146 1133
rect -112 957 -106 1133
rect -152 945 -106 957
rect 106 1133 152 1145
rect 106 957 112 1133
rect 146 957 152 1133
rect 106 945 152 957
rect -96 907 96 913
rect -96 873 -84 907
rect 84 873 96 907
rect -96 867 96 873
rect -96 799 96 805
rect -96 765 -84 799
rect 84 765 96 799
rect -96 759 96 765
rect -152 715 -106 727
rect -152 539 -146 715
rect -112 539 -106 715
rect -152 527 -106 539
rect 106 715 152 727
rect 106 539 112 715
rect 146 539 152 715
rect 106 527 152 539
rect -96 489 96 495
rect -96 455 -84 489
rect 84 455 96 489
rect -96 449 96 455
rect -96 381 96 387
rect -96 347 -84 381
rect 84 347 96 381
rect -96 341 96 347
rect -152 297 -106 309
rect -152 121 -146 297
rect -112 121 -106 297
rect -152 109 -106 121
rect 106 297 152 309
rect 106 121 112 297
rect 146 121 152 297
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -297 -146 -121
rect -112 -297 -106 -121
rect -152 -309 -106 -297
rect 106 -121 152 -109
rect 106 -297 112 -121
rect 146 -297 152 -121
rect 106 -309 152 -297
rect -96 -347 96 -341
rect -96 -381 -84 -347
rect 84 -381 96 -347
rect -96 -387 96 -381
rect -96 -455 96 -449
rect -96 -489 -84 -455
rect 84 -489 96 -455
rect -96 -495 96 -489
rect -152 -539 -106 -527
rect -152 -715 -146 -539
rect -112 -715 -106 -539
rect -152 -727 -106 -715
rect 106 -539 152 -527
rect 106 -715 112 -539
rect 146 -715 152 -539
rect 106 -727 152 -715
rect -96 -765 96 -759
rect -96 -799 -84 -765
rect 84 -799 96 -765
rect -96 -805 96 -799
rect -96 -873 96 -867
rect -96 -907 -84 -873
rect 84 -907 96 -873
rect -96 -913 96 -907
rect -152 -957 -106 -945
rect -152 -1133 -146 -957
rect -112 -1133 -106 -957
rect -152 -1145 -106 -1133
rect 106 -957 152 -945
rect 106 -1133 112 -957
rect 146 -1133 152 -957
rect 106 -1145 152 -1133
rect -96 -1183 96 -1177
rect -96 -1217 -84 -1183
rect 84 -1217 96 -1183
rect -96 -1223 96 -1217
rect -96 -1291 96 -1285
rect -96 -1325 -84 -1291
rect 84 -1325 96 -1291
rect -96 -1331 96 -1325
rect -152 -1375 -106 -1363
rect -152 -1551 -146 -1375
rect -112 -1551 -106 -1375
rect -152 -1563 -106 -1551
rect 106 -1375 152 -1363
rect 106 -1551 112 -1375
rect 146 -1551 152 -1375
rect 106 -1563 152 -1551
rect -96 -1601 96 -1595
rect -96 -1635 -84 -1601
rect 84 -1635 96 -1601
rect -96 -1641 96 -1635
rect -238 -1703 238 -1697
rect -238 -1737 -226 -1703
rect 226 -1737 238 -1703
rect -238 -1743 238 -1737
<< properties >>
string FIXED_BBOX -243 -1720 243 1720
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
