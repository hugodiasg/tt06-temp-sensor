VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_hugodg_temp_sensor
  CLASS BLOCK ;
  FOREIGN tt_um_hugodg_temp_sensor ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.000000 ;
    ANTENNADIFFAREA 49.667625 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 30.224998 ;
    ANTENNADIFFAREA 18.850000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.225000 ;
    ANTENNADIFFAREA 12.156000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 120.200 179.840 129.800 196.800 ;
      LAYER nwell ;
        RECT 130.935 179.835 136.265 195.965 ;
        RECT 137.535 175.635 145.865 195.765 ;
        RECT 143.410 168.625 147.110 168.760 ;
        RECT 129.645 161.795 147.110 168.625 ;
      LAYER pwell ;
        RECT 132.310 153.360 143.310 160.260 ;
        RECT 132.310 153.260 137.210 153.360 ;
        RECT 139.410 153.260 143.310 153.360 ;
        RECT 132.310 144.300 143.310 153.260 ;
      LAYER nwell ;
        RECT 143.410 143.660 147.110 161.795 ;
        RECT 129.610 136.860 147.110 143.660 ;
        RECT 125.200 124.000 126.400 125.200 ;
      LAYER pwell ;
        RECT 123.545 123.665 124.225 123.805 ;
        RECT 123.355 123.495 124.225 123.665 ;
        RECT 123.545 119.295 124.225 123.495 ;
      LAYER nwell ;
        RECT 124.745 123.100 126.400 124.000 ;
      LAYER pwell ;
        RECT 123.545 118.365 124.445 119.295 ;
        RECT 123.545 115.645 124.225 118.365 ;
        RECT 123.545 113.290 124.455 115.645 ;
      LAYER nwell ;
        RECT 124.745 113.040 126.350 123.100 ;
      LAYER pwell ;
        RECT 120.720 109.620 123.820 111.730 ;
      LAYER nwell ;
        RECT 124.070 109.620 129.260 111.730 ;
      LAYER pwell ;
        RECT 130.000 109.040 149.100 125.000 ;
      LAYER li1 ;
        RECT 120.380 196.450 129.620 196.620 ;
        RECT 120.380 195.700 120.550 196.450 ;
        RECT 121.470 195.770 122.510 195.940 ;
        RECT 123.560 195.770 124.600 195.940 ;
        RECT 125.650 195.770 126.690 195.940 ;
        RECT 127.740 195.770 128.780 195.940 ;
        RECT 120.380 194.600 120.600 195.700 ;
        RECT 121.130 194.710 121.300 195.710 ;
        RECT 122.680 194.710 122.850 195.710 ;
        RECT 123.220 194.710 123.390 195.710 ;
        RECT 124.770 194.710 124.940 195.710 ;
        RECT 125.310 194.710 125.480 195.710 ;
        RECT 126.860 194.710 127.030 195.710 ;
        RECT 127.400 194.710 127.570 195.710 ;
        RECT 128.950 194.710 129.120 195.710 ;
        RECT 120.380 191.300 120.550 194.600 ;
        RECT 121.470 194.480 122.510 194.650 ;
        RECT 123.560 194.480 124.600 194.650 ;
        RECT 125.650 194.480 126.690 194.650 ;
        RECT 127.740 194.480 128.780 194.650 ;
        RECT 121.470 193.870 122.510 194.040 ;
        RECT 123.560 193.870 124.600 194.040 ;
        RECT 125.650 193.870 126.690 194.040 ;
        RECT 127.740 193.870 128.780 194.040 ;
        RECT 121.130 192.810 121.300 193.810 ;
        RECT 122.680 192.810 122.850 193.810 ;
        RECT 123.220 192.810 123.390 193.810 ;
        RECT 124.770 192.810 124.940 193.810 ;
        RECT 125.310 192.810 125.480 193.810 ;
        RECT 126.860 192.810 127.030 193.810 ;
        RECT 127.400 192.810 127.570 193.810 ;
        RECT 128.950 192.810 129.120 193.810 ;
        RECT 121.470 192.580 122.510 192.750 ;
        RECT 123.560 192.580 124.600 192.750 ;
        RECT 125.650 192.580 126.690 192.750 ;
        RECT 127.740 192.580 128.780 192.750 ;
        RECT 121.470 191.970 122.510 192.140 ;
        RECT 123.560 191.970 124.600 192.140 ;
        RECT 125.650 191.970 126.690 192.140 ;
        RECT 127.740 191.970 128.780 192.140 ;
        RECT 120.380 190.200 120.600 191.300 ;
        RECT 121.130 190.910 121.300 191.910 ;
        RECT 122.680 190.910 122.850 191.910 ;
        RECT 123.220 190.910 123.390 191.910 ;
        RECT 124.770 190.910 124.940 191.910 ;
        RECT 125.310 190.910 125.480 191.910 ;
        RECT 126.860 190.910 127.030 191.910 ;
        RECT 127.400 190.910 127.570 191.910 ;
        RECT 128.950 190.910 129.120 191.910 ;
        RECT 121.470 190.680 122.510 190.850 ;
        RECT 123.560 190.680 124.600 190.850 ;
        RECT 125.650 190.680 126.690 190.850 ;
        RECT 127.740 190.680 128.780 190.850 ;
        RECT 120.380 186.700 120.550 190.200 ;
        RECT 121.470 190.070 122.510 190.240 ;
        RECT 123.560 190.070 124.600 190.240 ;
        RECT 125.650 190.070 126.690 190.240 ;
        RECT 127.740 190.070 128.780 190.240 ;
        RECT 121.130 189.010 121.300 190.010 ;
        RECT 122.680 189.010 122.850 190.010 ;
        RECT 123.220 189.010 123.390 190.010 ;
        RECT 124.770 189.010 124.940 190.010 ;
        RECT 125.310 189.010 125.480 190.010 ;
        RECT 126.860 189.010 127.030 190.010 ;
        RECT 127.400 189.010 127.570 190.010 ;
        RECT 128.950 189.010 129.120 190.010 ;
        RECT 121.470 188.780 122.510 188.950 ;
        RECT 123.560 188.780 124.600 188.950 ;
        RECT 125.650 188.780 126.690 188.950 ;
        RECT 127.740 188.780 128.780 188.950 ;
        RECT 121.470 188.170 122.510 188.340 ;
        RECT 123.560 188.170 124.600 188.340 ;
        RECT 125.650 188.170 126.690 188.340 ;
        RECT 127.740 188.170 128.780 188.340 ;
        RECT 121.130 187.110 121.300 188.110 ;
        RECT 122.680 187.110 122.850 188.110 ;
        RECT 123.220 187.110 123.390 188.110 ;
        RECT 124.770 187.110 124.940 188.110 ;
        RECT 125.310 187.110 125.480 188.110 ;
        RECT 126.860 187.110 127.030 188.110 ;
        RECT 127.400 187.110 127.570 188.110 ;
        RECT 128.950 187.110 129.120 188.110 ;
        RECT 121.470 186.880 122.510 187.050 ;
        RECT 123.560 186.880 124.600 187.050 ;
        RECT 125.650 186.880 126.690 187.050 ;
        RECT 127.740 186.880 128.780 187.050 ;
        RECT 120.380 185.600 120.600 186.700 ;
        RECT 121.470 186.270 122.510 186.440 ;
        RECT 123.560 186.270 124.600 186.440 ;
        RECT 125.650 186.270 126.690 186.440 ;
        RECT 127.740 186.270 128.780 186.440 ;
        RECT 120.380 182.500 120.550 185.600 ;
        RECT 121.130 185.210 121.300 186.210 ;
        RECT 122.680 185.210 122.850 186.210 ;
        RECT 123.220 185.210 123.390 186.210 ;
        RECT 124.770 185.210 124.940 186.210 ;
        RECT 125.310 185.210 125.480 186.210 ;
        RECT 126.860 185.210 127.030 186.210 ;
        RECT 127.400 185.210 127.570 186.210 ;
        RECT 128.950 185.210 129.120 186.210 ;
        RECT 121.470 184.980 122.510 185.150 ;
        RECT 123.560 184.980 124.600 185.150 ;
        RECT 125.650 184.980 126.690 185.150 ;
        RECT 127.740 184.980 128.780 185.150 ;
        RECT 121.470 184.370 122.510 184.540 ;
        RECT 123.560 184.370 124.600 184.540 ;
        RECT 125.650 184.370 126.690 184.540 ;
        RECT 127.740 184.370 128.780 184.540 ;
        RECT 121.130 183.310 121.300 184.310 ;
        RECT 122.680 183.310 122.850 184.310 ;
        RECT 123.220 183.310 123.390 184.310 ;
        RECT 124.770 183.310 124.940 184.310 ;
        RECT 125.310 183.310 125.480 184.310 ;
        RECT 126.860 183.310 127.030 184.310 ;
        RECT 127.400 183.310 127.570 184.310 ;
        RECT 128.950 183.310 129.120 184.310 ;
        RECT 121.470 183.080 122.510 183.250 ;
        RECT 123.560 183.080 124.600 183.250 ;
        RECT 125.650 183.080 126.690 183.250 ;
        RECT 127.740 183.080 128.780 183.250 ;
        RECT 120.380 181.400 120.600 182.500 ;
        RECT 121.470 182.470 122.510 182.640 ;
        RECT 123.560 182.470 124.600 182.640 ;
        RECT 125.650 182.470 126.690 182.640 ;
        RECT 127.740 182.470 128.780 182.640 ;
        RECT 121.130 181.410 121.300 182.410 ;
        RECT 122.680 181.410 122.850 182.410 ;
        RECT 123.220 181.410 123.390 182.410 ;
        RECT 124.770 181.410 124.940 182.410 ;
        RECT 125.310 181.410 125.480 182.410 ;
        RECT 126.860 181.410 127.030 182.410 ;
        RECT 127.400 181.410 127.570 182.410 ;
        RECT 128.950 181.410 129.120 182.410 ;
        RECT 120.380 180.190 120.550 181.400 ;
        RECT 121.470 181.180 122.510 181.350 ;
        RECT 123.560 181.180 124.600 181.350 ;
        RECT 125.650 181.180 126.690 181.350 ;
        RECT 127.740 181.180 128.780 181.350 ;
        RECT 129.450 180.190 129.620 196.450 ;
        RECT 120.380 180.020 129.620 180.190 ;
        RECT 131.115 195.615 136.085 195.785 ;
        RECT 131.115 180.185 131.285 195.615 ;
        RECT 132.680 194.790 134.720 194.960 ;
        RECT 132.295 193.730 132.465 194.730 ;
        RECT 134.935 193.730 135.105 194.730 ;
        RECT 132.680 193.500 134.720 193.670 ;
        RECT 132.680 192.890 134.720 193.060 ;
        RECT 132.295 191.830 132.465 192.830 ;
        RECT 134.935 191.830 135.105 192.830 ;
        RECT 132.680 191.600 134.720 191.770 ;
        RECT 132.295 190.540 132.465 191.540 ;
        RECT 134.935 190.540 135.105 191.540 ;
        RECT 132.680 190.310 134.720 190.480 ;
        RECT 132.295 189.250 132.465 190.250 ;
        RECT 134.935 189.250 135.105 190.250 ;
        RECT 132.680 189.020 134.720 189.190 ;
        RECT 132.295 187.960 132.465 188.960 ;
        RECT 134.935 187.960 135.105 188.960 ;
        RECT 132.680 187.730 134.720 187.900 ;
        RECT 132.295 186.670 132.465 187.670 ;
        RECT 134.935 186.670 135.105 187.670 ;
        RECT 132.680 186.440 134.720 186.610 ;
        RECT 132.295 185.380 132.465 186.380 ;
        RECT 134.935 185.380 135.105 186.380 ;
        RECT 132.680 185.150 134.720 185.320 ;
        RECT 132.295 184.090 132.465 185.090 ;
        RECT 134.935 184.090 135.105 185.090 ;
        RECT 132.680 183.860 134.720 184.030 ;
        RECT 132.295 182.800 132.465 183.800 ;
        RECT 134.935 182.800 135.105 183.800 ;
        RECT 132.680 182.570 134.720 182.740 ;
        RECT 132.680 181.990 134.720 182.160 ;
        RECT 132.295 180.930 132.465 181.930 ;
        RECT 134.935 180.930 135.105 181.930 ;
        RECT 132.680 180.700 134.720 180.870 ;
        RECT 134.100 180.185 134.600 180.400 ;
        RECT 135.915 180.185 136.085 195.615 ;
        RECT 131.115 180.015 136.085 180.185 ;
        RECT 137.715 195.415 145.685 195.585 ;
        RECT 134.100 180.000 134.600 180.015 ;
        RECT 137.715 175.985 137.885 195.415 ;
        RECT 138.880 194.690 140.920 194.860 ;
        RECT 138.495 193.630 138.665 194.630 ;
        RECT 141.135 193.630 141.305 194.630 ;
        RECT 138.880 193.400 140.920 193.570 ;
        RECT 138.880 192.790 140.920 192.960 ;
        RECT 138.495 191.730 138.665 192.730 ;
        RECT 141.135 191.730 141.305 192.730 ;
        RECT 145.515 192.600 145.685 195.415 ;
        RECT 145.500 191.800 145.700 192.600 ;
        RECT 138.880 191.500 140.920 191.670 ;
        RECT 138.495 190.440 138.665 191.440 ;
        RECT 141.135 190.440 141.305 191.440 ;
        RECT 138.880 190.210 140.920 190.380 ;
        RECT 138.880 189.590 140.920 189.760 ;
        RECT 138.495 188.530 138.665 189.530 ;
        RECT 141.135 188.530 141.305 189.530 ;
        RECT 138.880 188.300 140.920 188.470 ;
        RECT 138.495 187.240 138.665 188.240 ;
        RECT 141.135 187.240 141.305 188.240 ;
        RECT 142.280 187.790 144.320 187.960 ;
        RECT 138.880 187.010 140.920 187.180 ;
        RECT 138.495 185.950 138.665 186.950 ;
        RECT 141.135 185.950 141.305 186.950 ;
        RECT 141.895 186.730 142.065 187.730 ;
        RECT 144.535 186.730 144.705 187.730 ;
        RECT 145.515 187.000 145.685 191.800 ;
        RECT 142.280 186.500 144.320 186.670 ;
        RECT 145.500 186.200 145.700 187.000 ;
        RECT 142.280 185.890 144.320 186.060 ;
        RECT 138.880 185.720 140.920 185.890 ;
        RECT 138.495 184.660 138.665 185.660 ;
        RECT 141.135 184.660 141.305 185.660 ;
        RECT 141.895 184.830 142.065 185.830 ;
        RECT 144.535 184.830 144.705 185.830 ;
        RECT 142.280 184.600 144.320 184.770 ;
        RECT 138.880 184.430 140.920 184.600 ;
        RECT 142.280 183.990 144.320 184.160 ;
        RECT 138.880 183.790 140.920 183.960 ;
        RECT 138.495 182.730 138.665 183.730 ;
        RECT 141.135 182.730 141.305 183.730 ;
        RECT 138.880 182.500 140.920 182.670 ;
        RECT 138.495 181.440 138.665 182.440 ;
        RECT 141.135 181.440 141.305 182.440 ;
        RECT 138.880 181.210 140.920 181.380 ;
        RECT 138.495 180.150 138.665 181.150 ;
        RECT 141.135 180.150 141.305 181.150 ;
        RECT 138.880 179.920 140.920 180.090 ;
        RECT 138.495 178.860 138.665 179.860 ;
        RECT 141.135 178.860 141.305 179.860 ;
        RECT 141.895 178.930 142.065 183.930 ;
        RECT 144.535 178.930 144.705 183.930 ;
        RECT 145.515 183.100 145.685 186.200 ;
        RECT 145.500 182.300 145.700 183.100 ;
        RECT 138.880 178.630 140.920 178.800 ;
        RECT 142.280 178.700 144.320 178.870 ;
        RECT 145.515 178.500 145.685 182.300 ;
        RECT 138.880 177.990 140.920 178.160 ;
        RECT 142.280 178.090 144.320 178.260 ;
        RECT 138.495 176.930 138.665 177.930 ;
        RECT 141.135 176.930 141.305 177.930 ;
        RECT 141.895 177.030 142.065 178.030 ;
        RECT 144.535 177.030 144.705 178.030 ;
        RECT 145.500 177.700 145.700 178.500 ;
        RECT 138.880 176.700 140.920 176.870 ;
        RECT 142.280 176.800 144.320 176.970 ;
        RECT 145.515 175.985 145.685 177.700 ;
        RECT 137.715 175.815 145.685 175.985 ;
        RECT 129.825 168.275 146.895 168.445 ;
        RECT 129.825 162.145 129.995 168.275 ;
        RECT 143.625 168.260 143.795 168.275 ;
        RECT 130.790 167.750 145.830 167.920 ;
        RECT 130.405 166.690 130.575 167.690 ;
        RECT 146.045 166.690 146.215 167.690 ;
        RECT 130.790 166.460 145.830 166.630 ;
        RECT 130.405 165.400 130.575 166.400 ;
        RECT 146.045 165.400 146.215 166.400 ;
        RECT 130.790 165.170 145.830 165.340 ;
        RECT 130.405 164.110 130.575 165.110 ;
        RECT 146.045 164.110 146.215 165.110 ;
        RECT 130.790 163.880 145.830 164.050 ;
        RECT 130.405 162.820 130.575 163.820 ;
        RECT 146.045 162.820 146.215 163.820 ;
        RECT 130.790 162.590 145.830 162.760 ;
        RECT 143.225 162.145 143.795 162.160 ;
        RECT 129.825 162.060 143.795 162.145 ;
        RECT 129.825 161.975 143.810 162.060 ;
        RECT 143.610 160.760 143.810 161.975 ;
        RECT 144.790 161.950 145.830 162.120 ;
        RECT 144.405 160.890 144.575 161.890 ;
        RECT 146.045 160.890 146.215 161.890 ;
        RECT 146.725 161.445 146.895 168.275 ;
        RECT 146.710 161.275 146.895 161.445 ;
        RECT 132.490 159.910 143.230 160.080 ;
        RECT 132.490 156.260 132.660 159.910 ;
        RECT 137.830 158.530 138.870 158.700 ;
        RECT 137.490 157.470 137.660 158.470 ;
        RECT 139.040 157.470 139.210 158.470 ;
        RECT 137.830 157.240 138.870 157.410 ;
        RECT 132.410 155.760 132.810 156.260 ;
        RECT 137.490 156.180 137.660 157.180 ;
        RECT 139.040 156.180 139.210 157.180 ;
        RECT 137.830 155.950 138.870 156.120 ;
        RECT 132.490 149.160 132.660 155.760 ;
        RECT 137.490 154.890 137.660 155.890 ;
        RECT 139.040 154.890 139.210 155.890 ;
        RECT 137.830 154.660 138.870 154.830 ;
        RECT 137.490 153.600 137.660 154.600 ;
        RECT 139.040 153.600 139.210 154.600 ;
        RECT 137.830 153.370 138.870 153.540 ;
        RECT 140.590 153.110 140.760 153.440 ;
        RECT 140.930 153.430 142.470 153.600 ;
        RECT 140.930 152.950 142.470 153.120 ;
        RECT 133.530 152.730 138.570 152.900 ;
        RECT 133.190 151.670 133.360 152.670 ;
        RECT 138.740 151.670 138.910 152.670 ;
        RECT 140.590 152.150 140.760 152.480 ;
        RECT 140.930 152.470 142.470 152.640 ;
        RECT 142.640 152.630 142.810 152.960 ;
        RECT 140.930 151.990 142.470 152.160 ;
        RECT 133.530 151.440 138.570 151.610 ;
        RECT 140.930 151.510 142.470 151.680 ;
        RECT 142.640 151.670 142.810 152.000 ;
        RECT 133.190 150.380 133.360 151.380 ;
        RECT 138.740 150.380 138.910 151.380 ;
        RECT 133.530 150.150 138.570 150.320 ;
        RECT 132.410 148.660 132.810 149.160 ;
        RECT 133.190 149.090 133.360 150.090 ;
        RECT 138.740 149.090 138.910 150.090 ;
        RECT 133.530 148.860 138.570 149.030 ;
        RECT 132.490 144.650 132.660 148.660 ;
        RECT 133.190 147.800 133.360 148.800 ;
        RECT 138.740 147.800 138.910 148.800 ;
        RECT 133.530 147.570 138.570 147.740 ;
        RECT 133.190 146.510 133.360 147.510 ;
        RECT 138.740 146.510 138.910 147.510 ;
        RECT 133.530 146.280 138.570 146.450 ;
        RECT 133.190 145.220 133.360 146.220 ;
        RECT 138.740 145.220 138.910 146.220 ;
        RECT 133.530 144.990 138.570 145.160 ;
        RECT 143.060 144.650 143.230 159.910 ;
        RECT 132.490 144.480 143.230 144.650 ;
        RECT 143.625 143.445 143.795 160.760 ;
        RECT 144.790 160.660 145.830 160.830 ;
        RECT 144.405 159.600 144.575 160.600 ;
        RECT 146.045 159.600 146.215 160.600 ;
        RECT 144.790 159.370 145.830 159.540 ;
        RECT 144.405 158.310 144.575 159.310 ;
        RECT 146.045 158.310 146.215 159.310 ;
        RECT 144.790 158.080 145.830 158.250 ;
        RECT 144.405 157.020 144.575 158.020 ;
        RECT 146.045 157.020 146.215 158.020 ;
        RECT 144.790 156.790 145.830 156.960 ;
        RECT 144.405 155.730 144.575 156.730 ;
        RECT 146.045 155.730 146.215 156.730 ;
        RECT 144.790 155.500 145.830 155.670 ;
        RECT 144.405 154.440 144.575 155.440 ;
        RECT 146.045 154.440 146.215 155.440 ;
        RECT 146.725 155.360 146.895 161.275 ;
        RECT 144.790 154.210 145.830 154.380 ;
        RECT 144.405 153.150 144.575 154.150 ;
        RECT 146.045 153.150 146.215 154.150 ;
        RECT 144.790 152.920 145.830 153.090 ;
        RECT 144.790 152.350 145.830 152.520 ;
        RECT 144.405 151.270 144.575 152.290 ;
        RECT 146.045 151.290 146.215 152.290 ;
        RECT 144.790 151.060 145.830 151.230 ;
        RECT 144.405 149.980 144.575 151.000 ;
        RECT 146.045 150.000 146.215 151.000 ;
        RECT 146.710 150.160 146.910 155.360 ;
        RECT 144.790 149.770 145.830 149.940 ;
        RECT 144.405 148.690 144.575 149.710 ;
        RECT 146.045 148.710 146.215 149.710 ;
        RECT 144.790 148.480 145.830 148.650 ;
        RECT 144.405 147.400 144.575 148.420 ;
        RECT 146.045 147.420 146.215 148.420 ;
        RECT 144.790 147.190 145.830 147.360 ;
        RECT 144.405 146.110 144.575 147.130 ;
        RECT 146.045 146.130 146.215 147.130 ;
        RECT 144.790 145.900 145.830 146.070 ;
        RECT 144.405 144.840 144.575 145.840 ;
        RECT 146.045 144.840 146.215 145.840 ;
        RECT 144.790 144.610 145.830 144.780 ;
        RECT 144.405 143.530 144.575 144.550 ;
        RECT 146.045 143.550 146.215 144.550 ;
        RECT 146.725 143.945 146.895 150.160 ;
        RECT 146.710 143.775 146.895 143.945 ;
        RECT 129.825 143.275 143.810 143.445 ;
        RECT 144.790 143.320 145.830 143.490 ;
        RECT 129.825 137.245 129.995 143.275 ;
        RECT 130.790 142.750 145.830 142.920 ;
        RECT 130.405 141.690 130.575 142.690 ;
        RECT 146.045 141.690 146.215 142.690 ;
        RECT 130.790 141.460 145.830 141.630 ;
        RECT 130.405 140.400 130.575 141.400 ;
        RECT 146.045 140.400 146.215 141.400 ;
        RECT 130.790 140.170 145.830 140.340 ;
        RECT 130.405 139.110 130.575 140.110 ;
        RECT 146.045 139.110 146.215 140.110 ;
        RECT 130.790 138.880 145.830 139.050 ;
        RECT 130.405 137.820 130.575 138.820 ;
        RECT 146.045 137.820 146.215 138.820 ;
        RECT 130.790 137.590 145.830 137.760 ;
        RECT 146.725 137.560 146.895 143.775 ;
        RECT 143.625 137.245 143.795 137.260 ;
        RECT 146.710 137.245 146.910 137.560 ;
        RECT 129.825 137.075 146.910 137.245 ;
        RECT 146.710 137.060 146.910 137.075 ;
        RECT 125.500 124.200 125.950 124.700 ;
        RECT 130.180 124.650 148.920 124.820 ;
        RECT 123.355 123.295 123.525 123.810 ;
        RECT 123.785 123.465 124.245 123.720 ;
        RECT 123.355 122.965 123.905 123.295 ;
        RECT 124.075 123.200 124.245 123.465 ;
        RECT 124.415 123.370 125.065 123.720 ;
        RECT 125.235 123.465 125.905 123.720 ;
        RECT 125.235 123.200 125.405 123.465 ;
        RECT 126.075 123.295 126.245 123.810 ;
        RECT 124.075 122.970 125.405 123.200 ;
        RECT 125.575 122.965 126.245 123.295 ;
        RECT 123.355 122.265 123.525 122.965 ;
        RECT 123.785 122.625 125.905 122.795 ;
        RECT 125.105 122.395 125.890 122.455 ;
        RECT 123.355 121.935 123.885 122.265 ;
        RECT 124.055 122.130 125.890 122.395 ;
        RECT 124.055 121.935 125.105 122.130 ;
        RECT 126.075 121.960 126.245 122.965 ;
        RECT 123.355 119.335 123.525 121.935 ;
        RECT 123.745 121.595 125.445 121.765 ;
        RECT 125.615 121.710 126.245 121.960 ;
        RECT 123.745 121.270 123.915 121.595 ;
        RECT 125.275 121.540 125.445 121.595 ;
        RECT 124.205 121.075 124.825 121.425 ;
        RECT 125.275 121.370 125.905 121.540 ;
        RECT 125.575 121.290 125.905 121.370 ;
        RECT 123.745 120.380 123.915 121.065 ;
        RECT 125.015 120.905 125.405 121.200 ;
        RECT 124.205 120.735 125.405 120.905 ;
        RECT 124.205 120.550 124.425 120.735 ;
        RECT 125.575 120.565 125.905 121.075 ;
        RECT 124.625 120.395 125.905 120.565 ;
        RECT 124.625 120.380 124.795 120.395 ;
        RECT 123.745 120.210 124.795 120.380 ;
        RECT 123.355 119.005 123.985 119.335 ;
        RECT 124.205 119.215 124.455 120.005 ;
        RECT 124.625 119.045 124.795 120.210 ;
        RECT 125.305 120.055 125.815 120.225 ;
        RECT 123.355 117.105 123.525 119.005 ;
        RECT 124.445 118.875 124.795 119.045 ;
        RECT 123.715 118.705 124.275 118.795 ;
        RECT 124.965 118.705 125.135 120.035 ;
        RECT 125.305 119.320 125.475 120.055 ;
        RECT 126.075 119.820 126.245 121.710 ;
        RECT 125.645 119.490 126.245 119.820 ;
        RECT 125.305 119.150 125.815 119.320 ;
        RECT 126.075 118.855 126.245 119.490 ;
        RECT 123.715 118.535 125.445 118.705 ;
        RECT 123.715 118.445 123.885 118.535 ;
        RECT 123.695 117.445 123.975 118.225 ;
        RECT 124.145 118.135 125.105 118.345 ;
        RECT 125.275 118.315 125.445 118.535 ;
        RECT 125.615 118.485 126.245 118.855 ;
        RECT 125.275 118.145 125.905 118.315 ;
        RECT 124.145 117.615 124.765 117.965 ;
        RECT 124.935 117.840 125.105 118.135 ;
        RECT 124.935 117.670 125.395 117.840 ;
        RECT 123.695 117.275 124.925 117.445 ;
        RECT 125.095 117.380 125.395 117.670 ;
        RECT 124.755 117.210 124.925 117.275 ;
        RECT 125.565 117.210 125.905 117.910 ;
        RECT 123.355 116.915 123.965 117.105 ;
        RECT 123.355 115.475 123.525 116.915 ;
        RECT 124.135 116.885 124.585 117.105 ;
        RECT 124.755 117.040 125.905 117.210 ;
        RECT 124.135 116.745 124.305 116.885 ;
        RECT 123.735 116.575 124.305 116.745 ;
        RECT 123.735 115.995 123.905 116.575 ;
        RECT 124.475 116.405 124.845 116.705 ;
        RECT 124.075 116.165 124.845 116.405 ;
        RECT 123.735 115.820 124.735 115.995 ;
        RECT 125.015 115.990 125.185 117.040 ;
        RECT 126.075 116.870 126.245 118.485 ;
        RECT 125.615 116.620 126.245 116.870 ;
        RECT 125.355 116.280 125.815 116.450 ;
        RECT 125.355 115.820 125.525 116.280 ;
        RECT 126.075 116.100 126.245 116.620 ;
        RECT 123.735 115.675 125.525 115.820 ;
        RECT 124.260 115.670 125.525 115.675 ;
        RECT 124.435 115.650 125.525 115.670 ;
        RECT 123.355 115.305 124.210 115.475 ;
        RECT 124.435 115.375 124.765 115.650 ;
        RECT 125.695 115.380 126.245 116.100 ;
        RECT 123.355 114.050 123.525 115.305 ;
        RECT 124.895 115.135 125.905 115.210 ;
        RECT 123.715 114.805 125.905 115.135 ;
        RECT 123.900 114.800 124.200 114.805 ;
        RECT 123.785 114.365 125.865 114.615 ;
        RECT 124.435 114.285 125.865 114.365 ;
        RECT 123.355 113.880 124.120 114.050 ;
        RECT 123.355 113.230 123.525 113.880 ;
        RECT 124.435 113.755 124.765 114.285 ;
        RECT 126.075 114.050 126.245 115.380 ;
        RECT 124.935 113.880 126.245 114.050 ;
        RECT 123.705 113.585 124.235 113.630 ;
        RECT 124.885 113.585 125.765 113.630 ;
        RECT 123.705 113.375 125.765 113.585 ;
        RECT 124.500 113.350 124.700 113.375 ;
        RECT 126.075 113.230 126.245 113.880 ;
        RECT 130.180 116.700 130.350 124.650 ;
        RECT 131.000 123.450 133.160 123.800 ;
        RECT 135.160 123.450 137.320 123.800 ;
        RECT 139.340 123.700 141.500 124.050 ;
        RECT 146.000 123.700 148.160 124.050 ;
        RECT 131.000 122.620 133.160 122.970 ;
        RECT 135.160 122.620 137.320 122.970 ;
        RECT 139.340 122.870 141.500 123.220 ;
        RECT 146.000 122.870 148.160 123.220 ;
        RECT 131.000 121.790 133.160 122.140 ;
        RECT 135.160 121.790 137.320 122.140 ;
        RECT 139.340 122.040 141.500 122.390 ;
        RECT 146.000 122.040 148.160 122.390 ;
        RECT 131.000 120.960 133.160 121.310 ;
        RECT 135.160 120.960 137.320 121.310 ;
        RECT 139.340 121.210 141.500 121.560 ;
        RECT 146.000 121.210 148.160 121.560 ;
        RECT 131.000 120.130 133.160 120.480 ;
        RECT 135.160 120.130 137.320 120.480 ;
        RECT 139.340 120.380 141.500 120.730 ;
        RECT 146.000 120.380 148.160 120.730 ;
        RECT 131.000 119.300 133.160 119.650 ;
        RECT 135.160 119.300 137.320 119.650 ;
        RECT 139.340 119.550 141.500 119.900 ;
        RECT 146.000 119.550 148.160 119.900 ;
        RECT 131.000 118.470 133.160 118.820 ;
        RECT 135.160 118.470 137.320 118.820 ;
        RECT 139.340 118.720 141.500 119.070 ;
        RECT 146.000 118.720 148.160 119.070 ;
        RECT 131.000 117.640 133.160 117.990 ;
        RECT 135.160 117.640 137.320 117.990 ;
        RECT 139.340 117.890 141.500 118.240 ;
        RECT 146.000 117.890 148.160 118.240 ;
        RECT 130.180 116.100 130.400 116.700 ;
        RECT 139.340 116.330 141.500 116.680 ;
        RECT 146.000 116.330 148.160 116.680 ;
        RECT 120.900 111.380 123.640 111.550 ;
        RECT 120.900 109.970 121.070 111.380 ;
        RECT 121.410 110.510 121.580 110.840 ;
        RECT 121.750 110.810 122.790 110.980 ;
        RECT 121.750 110.370 122.790 110.540 ;
        RECT 122.960 110.510 123.130 110.840 ;
        RECT 121.800 109.970 122.600 110.000 ;
        RECT 123.470 109.970 123.640 111.380 ;
        RECT 120.900 109.800 123.640 109.970 ;
        RECT 124.250 111.380 129.080 111.550 ;
        RECT 124.250 109.970 124.420 111.380 ;
        RECT 124.760 110.510 124.930 110.840 ;
        RECT 125.145 110.810 128.185 110.980 ;
        RECT 125.145 110.370 128.185 110.540 ;
        RECT 128.400 110.510 128.570 110.840 ;
        RECT 125.300 109.970 128.100 110.000 ;
        RECT 128.910 109.970 129.080 111.380 ;
        RECT 124.250 109.800 129.080 109.970 ;
        RECT 130.180 109.390 130.350 116.100 ;
        RECT 139.340 115.500 141.500 115.850 ;
        RECT 146.000 115.500 148.160 115.850 ;
        RECT 139.340 114.670 141.500 115.020 ;
        RECT 146.000 114.670 148.160 115.020 ;
        RECT 139.340 113.840 141.500 114.190 ;
        RECT 146.000 113.840 148.160 114.190 ;
        RECT 139.340 113.010 141.500 113.360 ;
        RECT 146.000 113.010 148.160 113.360 ;
        RECT 139.340 112.180 141.500 112.530 ;
        RECT 146.000 112.180 148.160 112.530 ;
        RECT 139.340 111.350 141.500 111.700 ;
        RECT 146.000 111.350 148.160 111.700 ;
        RECT 139.340 110.520 141.500 110.870 ;
        RECT 146.000 110.520 148.160 110.870 ;
        RECT 148.750 109.390 148.920 124.650 ;
        RECT 130.180 109.220 148.920 109.390 ;
      LAYER mcon ;
        RECT 121.550 195.770 122.430 195.940 ;
        RECT 123.640 195.770 124.520 195.940 ;
        RECT 125.730 195.770 126.610 195.940 ;
        RECT 127.820 195.770 128.700 195.940 ;
        RECT 120.400 194.600 120.600 195.700 ;
        RECT 121.130 194.790 121.300 195.630 ;
        RECT 122.680 194.790 122.850 195.630 ;
        RECT 123.220 194.790 123.390 195.630 ;
        RECT 124.770 194.790 124.940 195.630 ;
        RECT 125.310 194.790 125.480 195.630 ;
        RECT 126.860 194.790 127.030 195.630 ;
        RECT 127.400 194.790 127.570 195.630 ;
        RECT 128.950 194.790 129.120 195.630 ;
        RECT 121.550 194.480 122.430 194.650 ;
        RECT 123.640 194.480 124.520 194.650 ;
        RECT 125.730 194.480 126.610 194.650 ;
        RECT 127.820 194.480 128.700 194.650 ;
        RECT 121.550 193.870 122.430 194.040 ;
        RECT 123.640 193.870 124.520 194.040 ;
        RECT 125.730 193.870 126.610 194.040 ;
        RECT 127.820 193.870 128.700 194.040 ;
        RECT 121.130 192.890 121.300 193.730 ;
        RECT 122.680 192.890 122.850 193.730 ;
        RECT 123.220 192.890 123.390 193.730 ;
        RECT 124.770 192.890 124.940 193.730 ;
        RECT 125.310 192.890 125.480 193.730 ;
        RECT 126.860 192.890 127.030 193.730 ;
        RECT 127.400 192.890 127.570 193.730 ;
        RECT 128.950 192.890 129.120 193.730 ;
        RECT 121.550 192.580 122.430 192.750 ;
        RECT 123.640 192.580 124.520 192.750 ;
        RECT 125.730 192.580 126.610 192.750 ;
        RECT 127.820 192.580 128.700 192.750 ;
        RECT 121.550 191.970 122.430 192.140 ;
        RECT 123.640 191.970 124.520 192.140 ;
        RECT 125.730 191.970 126.610 192.140 ;
        RECT 127.820 191.970 128.700 192.140 ;
        RECT 120.400 190.200 120.600 191.300 ;
        RECT 121.130 190.990 121.300 191.830 ;
        RECT 122.680 190.990 122.850 191.830 ;
        RECT 123.220 190.990 123.390 191.830 ;
        RECT 124.770 190.990 124.940 191.830 ;
        RECT 125.310 190.990 125.480 191.830 ;
        RECT 126.860 190.990 127.030 191.830 ;
        RECT 127.400 190.990 127.570 191.830 ;
        RECT 128.950 190.990 129.120 191.830 ;
        RECT 121.550 190.680 122.430 190.850 ;
        RECT 123.640 190.680 124.520 190.850 ;
        RECT 125.730 190.680 126.610 190.850 ;
        RECT 127.820 190.680 128.700 190.850 ;
        RECT 121.550 190.070 122.430 190.240 ;
        RECT 123.640 190.070 124.520 190.240 ;
        RECT 125.730 190.070 126.610 190.240 ;
        RECT 127.820 190.070 128.700 190.240 ;
        RECT 121.130 189.090 121.300 189.930 ;
        RECT 122.680 189.090 122.850 189.930 ;
        RECT 123.220 189.090 123.390 189.930 ;
        RECT 124.770 189.090 124.940 189.930 ;
        RECT 125.310 189.090 125.480 189.930 ;
        RECT 126.860 189.090 127.030 189.930 ;
        RECT 127.400 189.090 127.570 189.930 ;
        RECT 128.950 189.090 129.120 189.930 ;
        RECT 121.550 188.780 122.430 188.950 ;
        RECT 123.640 188.780 124.520 188.950 ;
        RECT 125.730 188.780 126.610 188.950 ;
        RECT 127.820 188.780 128.700 188.950 ;
        RECT 121.550 188.170 122.430 188.340 ;
        RECT 123.640 188.170 124.520 188.340 ;
        RECT 125.730 188.170 126.610 188.340 ;
        RECT 127.820 188.170 128.700 188.340 ;
        RECT 121.130 187.190 121.300 188.030 ;
        RECT 122.680 187.190 122.850 188.030 ;
        RECT 123.220 187.190 123.390 188.030 ;
        RECT 124.770 187.190 124.940 188.030 ;
        RECT 125.310 187.190 125.480 188.030 ;
        RECT 126.860 187.190 127.030 188.030 ;
        RECT 127.400 187.190 127.570 188.030 ;
        RECT 128.950 187.190 129.120 188.030 ;
        RECT 121.550 186.880 122.430 187.050 ;
        RECT 123.640 186.880 124.520 187.050 ;
        RECT 125.730 186.880 126.610 187.050 ;
        RECT 127.820 186.880 128.700 187.050 ;
        RECT 120.400 185.600 120.600 186.700 ;
        RECT 121.550 186.270 122.430 186.440 ;
        RECT 123.640 186.270 124.520 186.440 ;
        RECT 125.730 186.270 126.610 186.440 ;
        RECT 127.820 186.270 128.700 186.440 ;
        RECT 121.130 185.290 121.300 186.130 ;
        RECT 122.680 185.290 122.850 186.130 ;
        RECT 123.220 185.290 123.390 186.130 ;
        RECT 124.770 185.290 124.940 186.130 ;
        RECT 125.310 185.290 125.480 186.130 ;
        RECT 126.860 185.290 127.030 186.130 ;
        RECT 127.400 185.290 127.570 186.130 ;
        RECT 128.950 185.290 129.120 186.130 ;
        RECT 121.550 184.980 122.430 185.150 ;
        RECT 123.640 184.980 124.520 185.150 ;
        RECT 125.730 184.980 126.610 185.150 ;
        RECT 127.820 184.980 128.700 185.150 ;
        RECT 121.550 184.370 122.430 184.540 ;
        RECT 123.640 184.370 124.520 184.540 ;
        RECT 125.730 184.370 126.610 184.540 ;
        RECT 127.820 184.370 128.700 184.540 ;
        RECT 121.130 183.390 121.300 184.230 ;
        RECT 122.680 183.390 122.850 184.230 ;
        RECT 123.220 183.390 123.390 184.230 ;
        RECT 124.770 183.390 124.940 184.230 ;
        RECT 125.310 183.390 125.480 184.230 ;
        RECT 126.860 183.390 127.030 184.230 ;
        RECT 127.400 183.390 127.570 184.230 ;
        RECT 128.950 183.390 129.120 184.230 ;
        RECT 121.550 183.080 122.430 183.250 ;
        RECT 123.640 183.080 124.520 183.250 ;
        RECT 125.730 183.080 126.610 183.250 ;
        RECT 127.820 183.080 128.700 183.250 ;
        RECT 120.400 181.400 120.600 182.500 ;
        RECT 121.550 182.470 122.430 182.640 ;
        RECT 123.640 182.470 124.520 182.640 ;
        RECT 125.730 182.470 126.610 182.640 ;
        RECT 127.820 182.470 128.700 182.640 ;
        RECT 121.130 181.490 121.300 182.330 ;
        RECT 122.680 181.490 122.850 182.330 ;
        RECT 123.220 181.490 123.390 182.330 ;
        RECT 124.770 181.490 124.940 182.330 ;
        RECT 125.310 181.490 125.480 182.330 ;
        RECT 126.860 181.490 127.030 182.330 ;
        RECT 127.400 181.490 127.570 182.330 ;
        RECT 128.950 181.490 129.120 182.330 ;
        RECT 121.550 181.180 122.430 181.350 ;
        RECT 123.640 181.180 124.520 181.350 ;
        RECT 125.730 181.180 126.610 181.350 ;
        RECT 127.820 181.180 128.700 181.350 ;
        RECT 133.615 194.790 134.555 194.960 ;
        RECT 132.295 193.810 132.465 194.650 ;
        RECT 134.935 193.810 135.105 194.650 ;
        RECT 133.615 193.500 134.555 193.670 ;
        RECT 132.845 192.890 133.785 193.060 ;
        RECT 132.295 191.910 132.465 192.750 ;
        RECT 134.935 191.910 135.105 192.750 ;
        RECT 133.615 191.600 134.555 191.770 ;
        RECT 132.295 190.620 132.465 191.460 ;
        RECT 134.935 190.620 135.105 191.460 ;
        RECT 132.845 190.310 133.785 190.480 ;
        RECT 132.295 189.330 132.465 190.170 ;
        RECT 134.935 189.330 135.105 190.170 ;
        RECT 133.615 189.020 134.555 189.190 ;
        RECT 132.295 188.040 132.465 188.880 ;
        RECT 134.935 188.040 135.105 188.880 ;
        RECT 132.845 187.730 133.785 187.900 ;
        RECT 132.295 186.750 132.465 187.590 ;
        RECT 134.935 186.750 135.105 187.590 ;
        RECT 133.615 186.440 134.555 186.610 ;
        RECT 132.295 185.460 132.465 186.300 ;
        RECT 134.935 185.460 135.105 186.300 ;
        RECT 132.845 185.150 133.785 185.320 ;
        RECT 132.295 184.170 132.465 185.010 ;
        RECT 134.935 184.170 135.105 185.010 ;
        RECT 133.615 183.860 134.555 184.030 ;
        RECT 132.295 182.880 132.465 183.720 ;
        RECT 134.935 182.880 135.105 183.720 ;
        RECT 132.845 182.570 133.785 182.740 ;
        RECT 133.615 181.990 134.555 182.160 ;
        RECT 132.295 181.010 132.465 181.850 ;
        RECT 134.935 181.010 135.105 181.850 ;
        RECT 133.615 180.700 134.555 180.870 ;
        RECT 139.815 194.690 140.755 194.860 ;
        RECT 138.495 193.710 138.665 194.550 ;
        RECT 141.135 193.710 141.305 194.550 ;
        RECT 139.815 193.400 140.755 193.570 ;
        RECT 139.045 192.790 139.985 192.960 ;
        RECT 138.495 191.810 138.665 192.650 ;
        RECT 141.135 191.810 141.305 192.650 ;
        RECT 145.500 191.800 145.700 192.600 ;
        RECT 139.815 191.500 140.755 191.670 ;
        RECT 138.495 190.520 138.665 191.360 ;
        RECT 141.135 190.520 141.305 191.360 ;
        RECT 139.045 190.210 139.985 190.380 ;
        RECT 139.045 189.590 139.985 189.760 ;
        RECT 138.495 188.610 138.665 189.450 ;
        RECT 141.135 188.610 141.305 189.450 ;
        RECT 139.815 188.300 140.755 188.470 ;
        RECT 138.495 187.320 138.665 188.160 ;
        RECT 141.135 187.320 141.305 188.160 ;
        RECT 143.215 187.790 144.155 187.960 ;
        RECT 139.045 187.010 139.985 187.180 ;
        RECT 138.495 186.030 138.665 186.870 ;
        RECT 141.135 186.030 141.305 186.870 ;
        RECT 141.895 186.810 142.065 187.650 ;
        RECT 144.535 186.810 144.705 187.650 ;
        RECT 143.215 186.500 144.155 186.670 ;
        RECT 145.500 186.200 145.700 187.000 ;
        RECT 142.360 185.890 144.240 186.060 ;
        RECT 139.815 185.720 140.755 185.890 ;
        RECT 138.495 184.740 138.665 185.580 ;
        RECT 141.135 184.740 141.305 185.580 ;
        RECT 141.895 184.910 142.065 185.750 ;
        RECT 144.535 184.910 144.705 185.750 ;
        RECT 142.360 184.600 144.240 184.770 ;
        RECT 139.045 184.430 139.985 184.600 ;
        RECT 142.360 183.990 144.240 184.160 ;
        RECT 139.045 183.790 139.985 183.960 ;
        RECT 138.495 182.810 138.665 183.650 ;
        RECT 141.135 182.810 141.305 183.650 ;
        RECT 139.815 182.500 140.755 182.670 ;
        RECT 138.495 181.520 138.665 182.360 ;
        RECT 141.135 181.520 141.305 182.360 ;
        RECT 139.045 181.210 139.985 181.380 ;
        RECT 138.495 180.230 138.665 181.070 ;
        RECT 141.135 180.230 141.305 181.070 ;
        RECT 139.815 179.920 140.755 180.090 ;
        RECT 138.495 178.940 138.665 179.780 ;
        RECT 141.135 178.940 141.305 179.780 ;
        RECT 141.895 179.010 142.065 183.850 ;
        RECT 144.535 179.010 144.705 183.850 ;
        RECT 145.500 182.300 145.700 183.100 ;
        RECT 139.045 178.630 139.985 178.800 ;
        RECT 142.360 178.700 144.240 178.870 ;
        RECT 139.045 177.990 139.985 178.160 ;
        RECT 143.215 178.090 144.155 178.260 ;
        RECT 138.495 177.010 138.665 177.850 ;
        RECT 141.135 177.010 141.305 177.850 ;
        RECT 141.895 177.110 142.065 177.950 ;
        RECT 144.535 177.110 144.705 177.950 ;
        RECT 145.500 177.700 145.700 178.500 ;
        RECT 139.045 176.700 139.985 176.870 ;
        RECT 143.215 176.800 144.155 176.970 ;
        RECT 138.225 167.750 145.665 167.920 ;
        RECT 130.405 166.770 130.575 167.610 ;
        RECT 130.955 166.460 138.395 166.630 ;
        RECT 146.045 165.480 146.215 166.320 ;
        RECT 138.225 165.170 145.665 165.340 ;
        RECT 146.045 164.190 146.215 165.030 ;
        RECT 130.955 163.880 138.395 164.050 ;
        RECT 130.405 162.900 130.575 163.740 ;
        RECT 138.225 162.590 145.665 162.760 ;
        RECT 144.955 161.950 145.395 162.120 ;
        RECT 144.405 160.970 144.575 161.810 ;
        RECT 137.995 158.530 138.435 158.700 ;
        RECT 137.490 157.550 137.660 158.390 ;
        RECT 139.040 157.550 139.210 158.390 ;
        RECT 138.265 157.240 138.705 157.410 ;
        RECT 137.490 156.260 137.660 157.100 ;
        RECT 132.410 155.760 132.810 156.260 ;
        RECT 139.040 156.260 139.210 157.100 ;
        RECT 137.995 155.950 138.435 156.120 ;
        RECT 137.490 154.970 137.660 155.810 ;
        RECT 139.040 154.970 139.210 155.810 ;
        RECT 138.265 154.660 138.705 154.830 ;
        RECT 137.490 153.680 137.660 154.520 ;
        RECT 139.040 153.680 139.210 154.520 ;
        RECT 137.995 153.370 138.435 153.540 ;
        RECT 141.095 153.430 141.785 153.600 ;
        RECT 140.590 153.190 140.760 153.360 ;
        RECT 141.615 152.950 142.305 153.120 ;
        RECT 135.965 152.730 138.405 152.900 ;
        RECT 142.640 152.710 142.810 152.880 ;
        RECT 133.190 151.750 133.360 152.590 ;
        RECT 138.740 151.750 138.910 152.590 ;
        RECT 141.095 152.470 141.785 152.640 ;
        RECT 140.590 152.230 140.760 152.400 ;
        RECT 141.615 151.990 142.305 152.160 ;
        RECT 142.640 151.750 142.810 151.920 ;
        RECT 133.695 151.440 136.135 151.610 ;
        RECT 141.095 151.510 141.785 151.680 ;
        RECT 133.190 150.460 133.360 151.300 ;
        RECT 138.740 150.460 138.910 151.300 ;
        RECT 135.965 150.150 138.405 150.320 ;
        RECT 133.190 149.170 133.360 150.010 ;
        RECT 132.410 148.660 132.810 149.160 ;
        RECT 138.740 149.170 138.910 150.010 ;
        RECT 133.695 148.860 136.135 149.030 ;
        RECT 133.190 147.880 133.360 148.720 ;
        RECT 138.740 147.880 138.910 148.720 ;
        RECT 135.965 147.570 138.405 147.740 ;
        RECT 133.190 146.590 133.360 147.430 ;
        RECT 138.740 146.590 138.910 147.430 ;
        RECT 133.695 146.280 136.135 146.450 ;
        RECT 133.190 145.300 133.360 146.140 ;
        RECT 138.740 145.300 138.910 146.140 ;
        RECT 135.965 144.990 138.405 145.160 ;
        RECT 145.225 160.660 145.665 160.830 ;
        RECT 144.405 159.680 144.575 160.520 ;
        RECT 146.045 159.680 146.215 160.520 ;
        RECT 144.955 159.370 145.395 159.540 ;
        RECT 144.405 158.390 144.575 159.230 ;
        RECT 145.225 158.080 145.665 158.250 ;
        RECT 144.405 157.100 144.575 157.940 ;
        RECT 144.955 156.790 145.395 156.960 ;
        RECT 144.405 155.810 144.575 156.650 ;
        RECT 145.225 155.500 145.665 155.670 ;
        RECT 144.405 154.520 144.575 155.360 ;
        RECT 144.955 154.210 145.395 154.380 ;
        RECT 144.405 153.230 144.575 154.070 ;
        RECT 145.225 152.920 145.665 153.090 ;
        RECT 144.955 152.350 145.395 152.520 ;
        RECT 145.225 151.060 145.665 151.230 ;
        RECT 146.710 150.160 146.910 155.360 ;
        RECT 144.955 149.770 145.395 149.940 ;
        RECT 145.225 148.480 145.665 148.650 ;
        RECT 144.955 147.190 145.395 147.360 ;
        RECT 145.225 145.900 145.665 146.070 ;
        RECT 144.405 144.920 144.575 145.760 ;
        RECT 146.045 144.920 146.215 145.760 ;
        RECT 144.955 144.610 145.395 144.780 ;
        RECT 145.225 143.320 145.665 143.490 ;
        RECT 138.225 142.750 145.665 142.920 ;
        RECT 130.405 141.770 130.575 142.610 ;
        RECT 130.955 141.460 138.395 141.630 ;
        RECT 146.045 140.480 146.215 141.320 ;
        RECT 138.225 140.170 145.665 140.340 ;
        RECT 146.045 139.190 146.215 140.030 ;
        RECT 130.955 138.880 138.395 139.050 ;
        RECT 130.405 137.900 130.575 138.740 ;
        RECT 138.225 137.590 145.665 137.760 ;
        RECT 125.650 124.300 125.900 124.650 ;
        RECT 123.355 123.495 123.525 123.665 ;
        RECT 123.355 123.035 123.525 123.205 ;
        RECT 124.500 123.500 124.800 123.700 ;
        RECT 126.075 123.495 126.245 123.665 ;
        RECT 124.545 123.030 124.715 123.200 ;
        RECT 126.075 123.035 126.245 123.205 ;
        RECT 123.355 122.575 123.525 122.745 ;
        RECT 125.225 122.625 125.395 122.795 ;
        RECT 126.075 122.575 126.245 122.745 ;
        RECT 123.355 122.115 123.525 122.285 ;
        RECT 124.150 122.000 124.350 122.300 ;
        RECT 126.075 122.115 126.245 122.285 ;
        RECT 123.355 121.655 123.525 121.825 ;
        RECT 123.355 121.195 123.525 121.365 ;
        RECT 126.075 121.655 126.245 121.825 ;
        RECT 124.545 121.195 124.715 121.365 ;
        RECT 123.355 120.735 123.525 120.905 ;
        RECT 123.355 120.275 123.525 120.445 ;
        RECT 126.075 121.195 126.245 121.365 ;
        RECT 125.225 120.735 125.395 120.905 ;
        RECT 126.075 120.735 126.245 120.905 ;
        RECT 126.075 120.275 126.245 120.445 ;
        RECT 123.355 119.815 123.525 119.985 ;
        RECT 123.355 119.355 123.525 119.525 ;
        RECT 124.205 119.835 124.375 120.005 ;
        RECT 124.205 119.475 124.375 119.645 ;
        RECT 123.355 118.895 123.525 119.065 ;
        RECT 123.355 118.435 123.525 118.605 ;
        RECT 126.075 119.815 126.245 119.985 ;
        RECT 126.075 119.355 126.245 119.525 ;
        RECT 126.075 118.895 126.245 119.065 ;
        RECT 123.355 117.975 123.525 118.145 ;
        RECT 123.355 117.515 123.525 117.685 ;
        RECT 126.075 118.435 126.245 118.605 ;
        RECT 124.545 117.615 124.715 117.785 ;
        RECT 126.075 117.975 126.245 118.145 ;
        RECT 125.225 117.615 125.395 117.785 ;
        RECT 123.355 117.055 123.525 117.225 ;
        RECT 123.355 116.595 123.525 116.765 ;
        RECT 126.075 117.515 126.245 117.685 ;
        RECT 126.075 117.055 126.245 117.225 ;
        RECT 123.355 116.135 123.525 116.305 ;
        RECT 123.355 115.675 123.525 115.845 ;
        RECT 124.520 116.535 124.690 116.705 ;
        RECT 124.205 116.235 124.375 116.405 ;
        RECT 126.075 116.595 126.245 116.765 ;
        RECT 126.075 116.135 126.245 116.305 ;
        RECT 126.075 115.675 126.245 115.845 ;
        RECT 123.355 115.215 123.525 115.385 ;
        RECT 126.075 115.215 126.245 115.385 ;
        RECT 123.355 114.755 123.525 114.925 ;
        RECT 126.075 114.755 126.245 114.925 ;
        RECT 123.355 114.295 123.525 114.465 ;
        RECT 126.075 114.295 126.245 114.465 ;
        RECT 123.355 113.835 123.525 114.005 ;
        RECT 126.075 113.835 126.245 114.005 ;
        RECT 123.355 113.375 123.525 113.545 ;
        RECT 126.075 113.375 126.245 113.545 ;
        RECT 131.090 123.530 133.075 123.720 ;
        RECT 135.245 123.530 137.230 123.720 ;
        RECT 139.430 123.780 141.415 123.970 ;
        RECT 146.085 123.780 148.070 123.970 ;
        RECT 131.090 122.700 133.075 122.890 ;
        RECT 135.245 122.700 137.230 122.890 ;
        RECT 139.430 122.950 141.415 123.140 ;
        RECT 146.085 122.950 148.070 123.140 ;
        RECT 131.090 121.870 133.075 122.060 ;
        RECT 135.245 121.870 137.230 122.060 ;
        RECT 139.430 122.120 141.415 122.310 ;
        RECT 146.085 122.120 148.070 122.310 ;
        RECT 131.090 121.040 133.075 121.230 ;
        RECT 135.245 121.040 137.230 121.230 ;
        RECT 139.430 121.290 141.415 121.480 ;
        RECT 146.085 121.290 148.070 121.480 ;
        RECT 131.090 120.210 133.075 120.400 ;
        RECT 135.245 120.210 137.230 120.400 ;
        RECT 139.430 120.460 141.415 120.650 ;
        RECT 146.085 120.460 148.070 120.650 ;
        RECT 131.090 119.380 133.075 119.570 ;
        RECT 135.245 119.380 137.230 119.570 ;
        RECT 139.430 119.630 141.415 119.820 ;
        RECT 146.085 119.630 148.070 119.820 ;
        RECT 131.090 118.550 133.075 118.740 ;
        RECT 135.245 118.550 137.230 118.740 ;
        RECT 139.430 118.800 141.415 118.990 ;
        RECT 146.085 118.800 148.070 118.990 ;
        RECT 131.090 117.720 133.075 117.910 ;
        RECT 135.245 117.720 137.230 117.910 ;
        RECT 139.430 117.970 141.415 118.160 ;
        RECT 146.085 117.970 148.070 118.160 ;
        RECT 139.430 116.410 141.415 116.600 ;
        RECT 146.085 116.410 148.070 116.600 ;
        RECT 121.830 110.810 122.710 110.980 ;
        RECT 121.410 110.590 121.580 110.760 ;
        RECT 122.960 110.590 123.130 110.760 ;
        RECT 121.830 110.370 122.710 110.540 ;
        RECT 121.800 109.800 122.600 110.000 ;
        RECT 125.225 110.810 128.105 110.980 ;
        RECT 124.760 110.590 124.930 110.760 ;
        RECT 128.400 110.590 128.570 110.760 ;
        RECT 125.225 110.370 128.105 110.540 ;
        RECT 125.300 109.800 128.100 110.000 ;
        RECT 139.430 115.580 141.415 115.770 ;
        RECT 146.085 115.580 148.070 115.770 ;
        RECT 139.430 114.750 141.415 114.940 ;
        RECT 146.085 114.750 148.070 114.940 ;
        RECT 139.430 113.920 141.415 114.110 ;
        RECT 146.085 113.920 148.070 114.110 ;
        RECT 139.430 113.090 141.415 113.280 ;
        RECT 146.085 113.090 148.070 113.280 ;
        RECT 139.430 112.260 141.415 112.450 ;
        RECT 146.085 112.260 148.070 112.450 ;
        RECT 139.430 111.430 141.415 111.620 ;
        RECT 146.085 111.430 148.070 111.620 ;
        RECT 139.430 110.600 141.415 110.790 ;
        RECT 146.085 110.600 148.070 110.790 ;
      LAYER met1 ;
        RECT 109.620 196.510 110.620 197.110 ;
        RECT 107.920 175.010 108.420 175.060 ;
        RECT 107.920 175.000 108.520 175.010 ;
        RECT 106.500 174.010 108.520 175.000 ;
        RECT 106.500 174.000 108.420 174.010 ;
        RECT 107.920 173.960 108.420 174.000 ;
        RECT 107.900 172.010 108.600 172.050 ;
        RECT 106.520 171.010 108.620 172.010 ;
        RECT 107.900 170.950 108.600 171.010 ;
        RECT 106.520 130.410 108.620 131.410 ;
        RECT 106.520 128.310 107.520 128.510 ;
        RECT 106.520 127.510 108.520 128.310 ;
        RECT 107.920 126.710 108.520 126.760 ;
        RECT 106.520 125.910 108.520 126.710 ;
        RECT 106.520 125.710 107.520 125.910 ;
        RECT 107.920 125.860 108.520 125.910 ;
        RECT 106.520 125.310 107.520 125.410 ;
        RECT 106.520 124.410 108.620 125.310 ;
        RECT 107.520 124.310 108.620 124.410 ;
        RECT 109.220 116.310 111.420 196.510 ;
        RECT 119.400 194.400 129.250 196.000 ;
        RECT 134.100 194.990 134.600 195.000 ;
        RECT 133.555 194.900 134.615 194.990 ;
        RECT 133.555 194.760 135.200 194.900 ;
        RECT 140.500 194.890 140.900 195.250 ;
        RECT 119.400 191.360 120.450 194.400 ;
        RECT 121.550 194.070 122.450 194.150 ;
        RECT 123.650 194.070 124.550 194.150 ;
        RECT 125.650 194.070 126.650 194.150 ;
        RECT 127.850 194.070 128.750 194.150 ;
        RECT 121.490 193.840 122.490 194.070 ;
        RECT 123.580 193.840 124.580 194.070 ;
        RECT 125.650 193.840 126.670 194.070 ;
        RECT 127.760 193.840 128.760 194.070 ;
        RECT 121.100 192.830 121.330 193.790 ;
        RECT 121.550 193.750 122.450 193.840 ;
        RECT 122.650 193.500 122.880 193.790 ;
        RECT 123.190 193.500 123.420 193.790 ;
        RECT 123.650 193.750 124.550 193.840 ;
        RECT 122.650 193.000 123.420 193.500 ;
        RECT 122.650 192.830 122.880 193.000 ;
        RECT 123.190 192.830 123.420 193.000 ;
        RECT 124.740 193.500 124.970 193.790 ;
        RECT 125.280 193.500 125.510 193.790 ;
        RECT 125.650 193.750 126.650 193.840 ;
        RECT 124.740 193.000 125.510 193.500 ;
        RECT 124.740 192.830 124.970 193.000 ;
        RECT 125.280 192.830 125.510 193.000 ;
        RECT 126.830 193.500 127.060 193.790 ;
        RECT 127.370 193.500 127.600 193.790 ;
        RECT 127.850 193.750 128.750 193.840 ;
        RECT 129.000 193.790 129.200 193.800 ;
        RECT 126.830 193.000 127.600 193.500 ;
        RECT 126.830 192.830 127.060 193.000 ;
        RECT 127.370 192.830 127.600 193.000 ;
        RECT 128.920 192.830 129.200 193.790 ;
        RECT 121.490 192.550 122.490 192.780 ;
        RECT 123.580 192.750 124.580 192.780 ;
        RECT 125.670 192.750 126.670 192.780 ;
        RECT 127.760 192.750 128.760 192.780 ;
        RECT 123.550 192.550 124.580 192.750 ;
        RECT 125.650 192.550 126.670 192.750 ;
        RECT 127.750 192.550 128.760 192.750 ;
        RECT 121.550 192.170 122.450 192.550 ;
        RECT 123.550 192.170 124.550 192.550 ;
        RECT 125.650 192.170 126.650 192.550 ;
        RECT 127.750 192.170 128.750 192.550 ;
        RECT 121.490 191.940 122.490 192.170 ;
        RECT 123.550 191.950 124.580 192.170 ;
        RECT 125.650 191.950 126.670 192.170 ;
        RECT 127.750 191.950 128.760 192.170 ;
        RECT 123.580 191.940 124.580 191.950 ;
        RECT 125.670 191.940 126.670 191.950 ;
        RECT 127.760 191.940 128.760 191.950 ;
        RECT 129.000 191.890 129.200 192.830 ;
        RECT 119.400 190.140 120.630 191.360 ;
        RECT 121.100 190.930 121.330 191.890 ;
        RECT 122.650 191.700 122.880 191.890 ;
        RECT 123.190 191.700 123.420 191.890 ;
        RECT 122.650 191.200 123.420 191.700 ;
        RECT 121.550 190.880 122.450 190.950 ;
        RECT 122.650 190.930 122.880 191.200 ;
        RECT 123.190 190.930 123.420 191.200 ;
        RECT 124.740 191.700 124.970 191.890 ;
        RECT 125.280 191.700 125.510 191.890 ;
        RECT 126.830 191.700 127.060 191.890 ;
        RECT 127.370 191.700 127.600 191.890 ;
        RECT 124.740 191.200 125.510 191.700 ;
        RECT 126.800 191.200 127.600 191.700 ;
        RECT 123.650 190.880 124.550 190.950 ;
        RECT 124.740 190.930 124.970 191.200 ;
        RECT 125.280 190.930 125.510 191.200 ;
        RECT 125.750 190.880 126.650 190.950 ;
        RECT 126.830 190.930 127.060 191.200 ;
        RECT 127.370 190.930 127.600 191.200 ;
        RECT 127.850 190.880 128.750 190.950 ;
        RECT 128.920 190.930 129.200 191.890 ;
        RECT 121.490 190.650 122.490 190.880 ;
        RECT 123.580 190.650 124.580 190.880 ;
        RECT 125.670 190.650 126.670 190.880 ;
        RECT 127.760 190.650 128.760 190.880 ;
        RECT 121.550 190.550 122.450 190.650 ;
        RECT 123.650 190.550 124.550 190.650 ;
        RECT 125.750 190.550 126.650 190.650 ;
        RECT 127.850 190.550 128.750 190.650 ;
        RECT 121.550 190.270 122.350 190.350 ;
        RECT 123.650 190.270 124.450 190.350 ;
        RECT 125.750 190.270 126.550 190.350 ;
        RECT 127.850 190.270 128.650 190.350 ;
        RECT 119.400 186.760 120.450 190.140 ;
        RECT 121.490 190.040 122.490 190.270 ;
        RECT 123.580 190.040 124.580 190.270 ;
        RECT 125.670 190.040 126.670 190.270 ;
        RECT 127.760 190.040 128.760 190.270 ;
        RECT 121.100 189.030 121.330 189.990 ;
        RECT 121.550 189.950 122.350 190.040 ;
        RECT 122.650 189.800 122.880 189.990 ;
        RECT 123.190 189.800 123.420 189.990 ;
        RECT 123.650 189.950 124.450 190.040 ;
        RECT 122.650 189.300 123.420 189.800 ;
        RECT 122.650 189.030 122.880 189.300 ;
        RECT 123.190 189.030 123.420 189.300 ;
        RECT 124.740 189.800 124.970 189.990 ;
        RECT 125.280 189.800 125.510 189.990 ;
        RECT 125.750 189.950 126.550 190.040 ;
        RECT 126.830 189.800 127.060 189.990 ;
        RECT 127.370 189.800 127.600 189.990 ;
        RECT 127.850 189.950 128.650 190.040 ;
        RECT 129.000 189.990 129.200 190.930 ;
        RECT 130.600 190.550 131.000 194.150 ;
        RECT 132.265 193.750 132.495 194.710 ;
        RECT 134.100 193.700 135.200 194.760 ;
        RECT 139.755 194.660 140.900 194.890 ;
        RECT 133.555 193.600 135.200 193.700 ;
        RECT 138.465 193.650 138.695 194.610 ;
        RECT 140.500 194.600 140.900 194.660 ;
        RECT 145.900 195.200 146.400 195.250 ;
        RECT 141.105 194.600 141.335 194.610 ;
        RECT 140.500 193.650 141.335 194.600 ;
        RECT 140.500 193.600 141.300 193.650 ;
        RECT 133.555 193.470 134.615 193.600 ;
        RECT 132.200 193.090 133.400 193.100 ;
        RECT 132.200 192.860 133.845 193.090 ;
        RECT 132.200 190.510 133.400 192.860 ;
        RECT 134.100 191.800 134.600 193.470 ;
        RECT 139.755 193.370 140.900 193.600 ;
        RECT 138.600 192.990 139.500 193.000 ;
        RECT 134.905 191.850 135.135 192.810 ;
        RECT 138.600 192.760 140.045 192.990 ;
        RECT 138.600 192.710 139.500 192.760 ;
        RECT 138.465 192.700 139.500 192.710 ;
        RECT 133.555 191.570 134.615 191.800 ;
        RECT 124.740 189.300 125.510 189.800 ;
        RECT 126.800 189.300 127.600 189.800 ;
        RECT 124.740 189.030 124.970 189.300 ;
        RECT 125.280 189.030 125.510 189.300 ;
        RECT 126.830 189.030 127.060 189.300 ;
        RECT 127.370 189.030 127.600 189.300 ;
        RECT 128.920 189.030 129.200 189.990 ;
        RECT 121.490 188.900 122.490 188.980 ;
        RECT 123.580 188.900 124.580 188.980 ;
        RECT 125.670 188.900 126.670 188.980 ;
        RECT 127.760 188.900 128.760 188.980 ;
        RECT 121.450 188.750 122.490 188.900 ;
        RECT 123.550 188.750 124.580 188.900 ;
        RECT 125.650 188.750 126.670 188.900 ;
        RECT 127.750 188.750 128.760 188.900 ;
        RECT 121.450 188.370 122.450 188.750 ;
        RECT 123.550 188.370 124.550 188.750 ;
        RECT 125.650 188.370 126.650 188.750 ;
        RECT 127.750 188.370 128.750 188.750 ;
        RECT 121.450 188.200 122.490 188.370 ;
        RECT 123.550 188.200 124.580 188.370 ;
        RECT 125.650 188.200 126.670 188.370 ;
        RECT 127.750 188.200 128.760 188.370 ;
        RECT 121.490 188.140 122.490 188.200 ;
        RECT 123.580 188.140 124.580 188.200 ;
        RECT 125.670 188.140 126.670 188.200 ;
        RECT 127.760 188.140 128.760 188.200 ;
        RECT 129.000 188.090 129.200 189.030 ;
        RECT 121.100 187.130 121.330 188.090 ;
        RECT 122.650 187.800 122.880 188.090 ;
        RECT 123.190 187.800 123.420 188.090 ;
        RECT 122.650 187.300 123.420 187.800 ;
        RECT 121.500 187.080 122.400 187.250 ;
        RECT 122.650 187.130 122.880 187.300 ;
        RECT 123.190 187.130 123.420 187.300 ;
        RECT 124.740 187.800 124.970 188.090 ;
        RECT 125.280 187.800 125.510 188.090 ;
        RECT 126.830 187.800 127.060 188.090 ;
        RECT 127.370 187.800 127.600 188.090 ;
        RECT 124.740 187.300 125.510 187.800 ;
        RECT 126.800 187.300 127.600 187.800 ;
        RECT 123.600 187.080 124.500 187.250 ;
        RECT 124.740 187.130 124.970 187.300 ;
        RECT 125.280 187.130 125.510 187.300 ;
        RECT 125.700 187.080 126.600 187.250 ;
        RECT 126.830 187.130 127.060 187.300 ;
        RECT 127.370 187.130 127.600 187.300 ;
        RECT 127.800 187.080 128.700 187.250 ;
        RECT 128.920 187.130 129.200 188.090 ;
        RECT 121.490 186.850 122.490 187.080 ;
        RECT 123.580 186.850 124.580 187.080 ;
        RECT 125.670 186.850 126.670 187.080 ;
        RECT 127.760 186.850 128.760 187.080 ;
        RECT 119.400 185.540 120.630 186.760 ;
        RECT 121.550 186.470 122.450 186.550 ;
        RECT 123.650 186.470 124.550 186.550 ;
        RECT 125.650 186.470 126.650 186.550 ;
        RECT 127.750 186.470 128.750 186.650 ;
        RECT 121.490 186.240 122.490 186.470 ;
        RECT 123.580 186.240 124.580 186.470 ;
        RECT 125.650 186.240 126.670 186.470 ;
        RECT 127.750 186.240 128.760 186.470 ;
        RECT 119.400 182.700 120.450 185.540 ;
        RECT 121.100 185.230 121.330 186.190 ;
        RECT 121.550 186.150 122.450 186.240 ;
        RECT 122.650 185.900 122.880 186.190 ;
        RECT 123.190 185.900 123.420 186.190 ;
        RECT 123.650 186.150 124.550 186.240 ;
        RECT 122.650 185.400 123.420 185.900 ;
        RECT 122.650 185.230 122.880 185.400 ;
        RECT 123.190 185.230 123.420 185.400 ;
        RECT 124.740 185.900 124.970 186.190 ;
        RECT 125.280 185.900 125.510 186.190 ;
        RECT 125.650 186.050 126.650 186.240 ;
        RECT 126.830 185.900 127.060 186.190 ;
        RECT 127.370 185.900 127.600 186.190 ;
        RECT 127.750 186.150 128.750 186.240 ;
        RECT 129.000 186.190 129.200 187.130 ;
        RECT 124.740 185.400 125.510 185.900 ;
        RECT 126.800 185.400 127.600 185.900 ;
        RECT 124.740 185.230 124.970 185.400 ;
        RECT 125.280 185.230 125.510 185.400 ;
        RECT 126.830 185.230 127.060 185.400 ;
        RECT 127.370 185.230 127.600 185.400 ;
        RECT 128.920 185.230 129.200 186.190 ;
        RECT 121.490 184.950 122.490 185.180 ;
        RECT 123.580 184.950 124.580 185.180 ;
        RECT 125.670 184.950 126.670 185.180 ;
        RECT 127.760 184.950 128.760 185.180 ;
        RECT 121.550 184.570 122.450 184.950 ;
        RECT 123.650 184.570 124.550 184.950 ;
        RECT 125.750 184.570 126.650 184.950 ;
        RECT 127.850 184.570 128.750 184.950 ;
        RECT 121.490 184.340 122.490 184.570 ;
        RECT 123.580 184.340 124.580 184.570 ;
        RECT 125.670 184.340 126.670 184.570 ;
        RECT 127.760 184.340 128.760 184.570 ;
        RECT 129.000 184.290 129.200 185.230 ;
        RECT 121.100 183.330 121.330 184.290 ;
        RECT 122.650 184.100 122.880 184.290 ;
        RECT 123.190 184.100 123.420 184.290 ;
        RECT 122.650 183.600 123.420 184.100 ;
        RECT 121.550 183.280 122.450 183.350 ;
        RECT 122.650 183.330 122.880 183.600 ;
        RECT 123.190 183.330 123.420 183.600 ;
        RECT 124.740 184.100 124.970 184.290 ;
        RECT 125.280 184.100 125.510 184.290 ;
        RECT 126.830 184.100 127.060 184.290 ;
        RECT 127.370 184.100 127.600 184.290 ;
        RECT 124.740 183.600 125.510 184.100 ;
        RECT 126.800 183.600 127.600 184.100 ;
        RECT 123.650 183.280 124.550 183.350 ;
        RECT 124.740 183.330 124.970 183.600 ;
        RECT 125.280 183.330 125.510 183.600 ;
        RECT 125.750 183.280 126.650 183.350 ;
        RECT 126.830 183.330 127.060 183.600 ;
        RECT 127.370 183.330 127.600 183.600 ;
        RECT 128.920 183.450 129.200 184.290 ;
        RECT 127.750 183.280 128.650 183.450 ;
        RECT 128.920 183.330 129.300 183.450 ;
        RECT 121.490 183.050 122.490 183.280 ;
        RECT 123.580 183.050 124.580 183.280 ;
        RECT 125.670 183.050 126.670 183.280 ;
        RECT 127.750 183.050 128.760 183.280 ;
        RECT 121.550 182.950 122.450 183.050 ;
        RECT 123.650 182.950 124.550 183.050 ;
        RECT 125.750 182.950 126.650 183.050 ;
        RECT 129.000 182.950 129.300 183.330 ;
        RECT 119.400 182.500 128.900 182.700 ;
        RECT 119.400 182.390 129.100 182.500 ;
        RECT 119.400 181.100 129.150 182.390 ;
        RECT 129.800 181.750 130.200 183.350 ;
        RECT 130.800 183.150 131.200 190.350 ;
        RECT 132.200 190.280 133.845 190.510 ;
        RECT 132.200 187.930 133.400 190.280 ;
        RECT 134.100 189.220 134.600 191.570 ;
        RECT 134.905 190.560 135.135 191.520 ;
        RECT 138.400 190.410 139.500 192.700 ;
        RECT 140.500 191.700 140.900 193.370 ;
        RECT 141.105 191.750 141.335 192.710 ;
        RECT 145.470 192.600 145.730 192.660 ;
        RECT 145.900 192.600 146.900 195.200 ;
        RECT 145.470 191.800 146.900 192.600 ;
        RECT 145.470 191.740 145.730 191.800 ;
        RECT 139.755 191.500 140.900 191.700 ;
        RECT 139.755 191.470 140.815 191.500 ;
        RECT 141.105 190.460 141.335 191.420 ;
        RECT 134.905 189.270 135.135 190.230 ;
        RECT 138.400 190.200 140.045 190.410 ;
        RECT 133.555 188.990 134.615 189.220 ;
        RECT 132.200 187.700 133.845 187.930 ;
        RECT 131.500 181.650 131.800 186.650 ;
        RECT 132.200 185.350 133.400 187.700 ;
        RECT 134.100 186.640 134.600 188.990 ;
        RECT 134.905 187.980 135.135 188.940 ;
        RECT 134.905 186.690 135.135 187.650 ;
        RECT 133.555 186.410 134.615 186.640 ;
        RECT 132.200 185.120 133.845 185.350 ;
        RECT 132.200 182.770 133.400 185.120 ;
        RECT 134.100 184.060 134.600 186.410 ;
        RECT 134.905 185.400 135.135 186.360 ;
        RECT 134.905 184.110 135.135 185.070 ;
        RECT 138.400 184.700 138.700 190.200 ;
        RECT 138.985 190.180 140.045 190.200 ;
        RECT 138.900 189.790 139.400 189.800 ;
        RECT 138.900 189.560 140.045 189.790 ;
        RECT 138.900 187.210 139.400 189.560 ;
        RECT 141.105 188.550 141.335 189.510 ;
        RECT 139.755 188.270 140.900 188.500 ;
        RECT 138.900 186.980 140.045 187.210 ;
        RECT 138.465 184.680 138.695 184.700 ;
        RECT 138.900 184.630 139.400 186.980 ;
        RECT 140.400 185.920 140.900 188.270 ;
        RECT 141.105 187.260 141.335 188.220 ;
        RECT 143.600 187.990 144.200 188.850 ;
        RECT 143.155 187.800 144.215 187.990 ;
        RECT 143.155 187.760 144.700 187.800 ;
        RECT 143.600 187.710 144.700 187.760 ;
        RECT 141.105 185.970 141.335 186.930 ;
        RECT 141.865 186.750 142.095 187.710 ;
        RECT 143.600 187.700 144.735 187.710 ;
        RECT 143.600 186.700 144.800 187.700 ;
        RECT 143.155 186.600 144.800 186.700 ;
        RECT 145.470 187.000 145.730 187.060 ;
        RECT 145.900 187.000 146.900 191.800 ;
        RECT 143.155 186.470 144.215 186.600 ;
        RECT 143.600 186.090 144.200 186.470 ;
        RECT 145.470 186.200 146.900 187.000 ;
        RECT 145.470 186.140 145.730 186.200 ;
        RECT 139.755 185.690 140.900 185.920 ;
        RECT 142.300 185.860 144.300 186.090 ;
        RECT 138.900 184.400 140.045 184.630 ;
        RECT 133.555 183.830 134.615 184.060 ;
        RECT 138.900 183.990 139.400 184.400 ;
        RECT 140.400 184.300 140.900 185.690 ;
        RECT 141.865 185.800 142.095 185.810 ;
        RECT 143.600 185.800 144.200 185.860 ;
        RECT 141.105 184.680 141.335 185.640 ;
        RECT 141.865 184.850 142.100 185.800 ;
        RECT 132.200 182.600 133.845 182.770 ;
        RECT 132.785 182.540 133.845 182.600 ;
        RECT 134.100 182.190 134.600 183.830 ;
        RECT 134.905 182.820 135.135 183.780 ;
        RECT 138.900 183.760 140.045 183.990 ;
        RECT 141.900 183.910 142.100 184.850 ;
        RECT 142.300 184.800 143.400 185.050 ;
        RECT 144.505 184.850 144.735 185.810 ;
        RECT 142.300 184.570 144.300 184.800 ;
        RECT 142.300 184.550 143.400 184.570 ;
        RECT 142.500 184.190 143.200 184.200 ;
        RECT 142.300 183.960 144.300 184.190 ;
        RECT 136.500 183.700 137.100 183.750 ;
        RECT 133.555 182.000 134.615 182.190 ;
        RECT 133.555 181.960 135.200 182.000 ;
        RECT 132.265 180.950 132.495 181.910 ;
        RECT 134.100 180.900 135.200 181.960 ;
        RECT 133.555 180.670 134.615 180.900 ;
        RECT 134.100 180.430 134.600 180.670 ;
        RECT 134.040 179.970 134.660 180.430 ;
        RECT 134.100 176.600 134.600 179.970 ;
        RECT 136.400 176.600 137.100 183.700 ;
        RECT 138.400 183.150 138.700 183.750 ;
        RECT 138.465 182.750 138.700 183.150 ;
        RECT 138.500 182.420 138.700 182.750 ;
        RECT 138.465 181.460 138.700 182.420 ;
        RECT 138.500 181.130 138.700 181.460 ;
        RECT 138.465 180.170 138.700 181.130 ;
        RECT 138.500 179.840 138.700 180.170 ;
        RECT 138.465 178.900 138.700 179.840 ;
        RECT 138.900 181.410 139.400 183.760 ;
        RECT 141.865 183.750 142.100 183.910 ;
        RECT 141.105 182.750 141.335 183.710 ;
        RECT 141.800 183.150 142.100 183.750 ;
        RECT 139.755 182.470 140.815 182.700 ;
        RECT 138.900 181.180 140.045 181.410 ;
        RECT 138.465 178.880 138.695 178.900 ;
        RECT 138.900 178.830 139.400 181.180 ;
        RECT 140.300 180.120 140.800 182.470 ;
        RECT 141.105 181.460 141.335 182.420 ;
        RECT 141.105 180.170 141.335 181.130 ;
        RECT 139.755 179.890 140.815 180.120 ;
        RECT 141.105 178.880 141.335 179.840 ;
        RECT 141.865 178.950 142.095 183.150 ;
        RECT 142.500 179.900 143.200 183.960 ;
        RECT 142.500 179.850 143.100 179.900 ;
        RECT 144.505 178.950 144.735 183.910 ;
        RECT 145.470 183.100 145.730 183.160 ;
        RECT 145.900 183.100 146.900 186.200 ;
        RECT 145.470 182.300 146.900 183.100 ;
        RECT 145.470 182.240 145.730 182.300 ;
        RECT 138.900 178.600 140.045 178.830 ;
        RECT 142.300 178.670 144.300 178.900 ;
        RECT 138.900 178.190 139.400 178.600 ;
        RECT 143.500 178.290 144.200 178.670 ;
        RECT 145.470 178.500 145.730 178.560 ;
        RECT 145.900 178.500 146.900 182.300 ;
        RECT 143.155 178.200 144.215 178.290 ;
        RECT 138.900 177.960 140.045 178.190 ;
        RECT 143.155 178.060 144.600 178.200 ;
        RECT 143.500 178.010 144.600 178.060 ;
        RECT 138.465 177.900 138.695 177.910 ;
        RECT 138.900 177.900 139.400 177.960 ;
        RECT 138.465 177.000 139.400 177.900 ;
        RECT 138.465 176.950 138.695 177.000 ;
        RECT 138.900 176.900 139.400 177.000 ;
        RECT 141.105 176.950 141.335 177.910 ;
        RECT 141.865 177.050 142.095 178.010 ;
        RECT 143.500 177.050 144.735 178.010 ;
        RECT 145.470 177.700 146.900 178.500 ;
        RECT 145.470 177.640 145.730 177.700 ;
        RECT 143.500 177.000 144.700 177.050 ;
        RECT 143.155 176.900 144.700 177.000 ;
        RECT 138.900 176.670 140.045 176.900 ;
        RECT 143.155 176.770 144.215 176.900 ;
        RECT 143.500 176.700 144.200 176.770 ;
        RECT 138.900 176.600 139.400 176.670 ;
        RECT 127.500 169.960 128.500 171.900 ;
        RECT 127.500 169.000 128.510 169.960 ;
        RECT 127.510 168.960 128.510 169.000 ;
        RECT 129.110 168.960 130.110 169.960 ;
        RECT 133.900 169.000 134.900 176.600 ;
        RECT 136.200 174.950 137.200 176.600 ;
        RECT 143.600 176.050 144.200 176.700 ;
        RECT 145.900 175.600 146.900 177.700 ;
        RECT 127.710 156.810 128.310 168.960 ;
        RECT 129.510 161.210 129.910 168.960 ;
        RECT 137.810 167.950 138.710 167.960 ;
        RECT 137.810 167.720 145.725 167.950 ;
        RECT 130.375 167.660 130.605 167.670 ;
        RECT 130.375 166.710 130.610 167.660 ;
        RECT 130.410 166.660 130.610 166.710 ;
        RECT 137.810 166.660 138.710 167.720 ;
        RECT 130.410 166.560 138.710 166.660 ;
        RECT 130.410 166.430 138.455 166.560 ;
        RECT 130.410 166.360 132.110 166.430 ;
        RECT 130.410 164.060 130.610 166.360 ;
        RECT 134.610 164.080 135.110 166.430 ;
        RECT 146.010 166.380 146.210 167.660 ;
        RECT 143.810 165.370 145.010 165.510 ;
        RECT 146.010 165.420 146.245 166.380 ;
        RECT 138.165 165.140 145.725 165.370 ;
        RECT 143.810 164.910 145.010 165.140 ;
        RECT 146.010 165.090 146.210 165.420 ;
        RECT 146.010 164.130 146.245 165.090 ;
        RECT 130.895 164.060 138.455 164.080 ;
        RECT 130.410 163.850 138.710 164.060 ;
        RECT 130.410 163.800 132.110 163.850 ;
        RECT 130.375 163.760 132.110 163.800 ;
        RECT 130.375 162.860 130.610 163.760 ;
        RECT 130.375 162.840 130.605 162.860 ;
        RECT 132.380 155.700 132.840 156.320 ;
        RECT 133.310 152.650 134.110 152.660 ;
        RECT 133.160 151.690 134.110 152.650 ;
        RECT 134.610 152.110 135.110 163.850 ;
        RECT 137.810 162.790 138.710 163.850 ;
        RECT 137.810 162.660 145.725 162.790 ;
        RECT 138.165 162.560 145.725 162.660 ;
        RECT 144.895 162.060 145.455 162.150 ;
        RECT 144.410 161.870 145.610 162.060 ;
        RECT 138.110 158.730 138.510 158.760 ;
        RECT 137.935 158.500 138.510 158.730 ;
        RECT 137.460 158.360 137.690 158.450 ;
        RECT 138.110 158.360 138.510 158.500 ;
        RECT 139.010 158.360 139.240 158.450 ;
        RECT 137.460 157.660 139.240 158.360 ;
        RECT 137.460 157.490 137.690 157.660 ;
        RECT 138.110 157.440 138.510 157.660 ;
        RECT 139.010 157.490 139.240 157.660 ;
        RECT 138.110 157.260 138.765 157.440 ;
        RECT 137.510 157.210 138.765 157.260 ;
        RECT 137.510 157.160 138.510 157.210 ;
        RECT 137.460 156.860 138.510 157.160 ;
        RECT 137.460 156.200 137.710 156.860 ;
        RECT 138.110 156.810 138.510 156.860 ;
        RECT 137.510 155.870 137.710 156.200 ;
        RECT 137.460 154.910 137.710 155.870 ;
        RECT 137.910 156.150 138.410 156.310 ;
        RECT 139.010 156.200 139.240 157.160 ;
        RECT 137.910 155.920 138.495 156.150 ;
        RECT 137.910 155.710 138.410 155.920 ;
        RECT 139.010 154.910 139.240 155.870 ;
        RECT 137.510 154.860 137.710 154.910 ;
        RECT 138.210 154.860 138.710 154.910 ;
        RECT 138.205 154.760 138.765 154.860 ;
        RECT 137.460 154.460 137.690 154.580 ;
        RECT 138.110 154.460 138.810 154.760 ;
        RECT 139.010 154.460 139.240 154.580 ;
        RECT 137.460 153.620 139.240 154.460 ;
        RECT 137.510 153.460 139.210 153.620 ;
        RECT 137.935 153.340 138.495 153.460 ;
        RECT 135.610 152.930 136.210 152.960 ;
        RECT 135.610 152.860 138.465 152.930 ;
        RECT 135.610 152.700 138.910 152.860 ;
        RECT 133.310 151.640 134.110 151.690 ;
        RECT 135.610 151.640 136.210 152.700 ;
        RECT 138.210 152.650 138.910 152.700 ;
        RECT 133.310 151.560 136.210 151.640 ;
        RECT 133.635 151.460 136.210 151.560 ;
        RECT 133.635 151.410 136.195 151.460 ;
        RECT 133.160 150.400 133.390 151.360 ;
        RECT 132.380 148.600 132.840 149.220 ;
        RECT 133.160 149.110 133.390 150.070 ;
        RECT 134.510 149.210 135.010 151.410 ;
        RECT 137.410 151.260 137.910 152.560 ;
        RECT 138.210 151.760 138.940 152.650 ;
        RECT 139.410 152.410 139.710 154.910 ;
        RECT 138.710 151.690 138.940 151.760 ;
        RECT 138.710 151.260 138.940 151.360 ;
        RECT 137.410 150.350 139.010 151.260 ;
        RECT 139.910 150.860 140.210 161.610 ;
        RECT 144.375 160.910 145.610 161.870 ;
        RECT 144.410 160.860 145.610 160.910 ;
        RECT 144.410 160.760 145.810 160.860 ;
        RECT 145.165 160.630 145.810 160.760 ;
        RECT 144.375 160.560 144.605 160.580 ;
        RECT 144.375 159.620 144.610 160.560 ;
        RECT 144.410 159.290 144.610 159.620 ;
        RECT 144.375 158.330 144.610 159.290 ;
        RECT 144.410 158.000 144.610 158.330 ;
        RECT 144.375 157.040 144.610 158.000 ;
        RECT 144.410 156.710 144.610 157.040 ;
        RECT 144.375 155.750 144.610 156.710 ;
        RECT 144.410 155.460 144.610 155.750 ;
        RECT 144.810 159.570 145.010 159.660 ;
        RECT 144.810 159.340 145.455 159.570 ;
        RECT 144.810 156.990 145.010 159.340 ;
        RECT 145.610 158.280 145.810 160.630 ;
        RECT 146.010 160.580 146.210 164.130 ;
        RECT 146.010 159.660 146.245 160.580 ;
        RECT 146.015 159.620 146.245 159.660 ;
        RECT 145.165 158.050 145.810 158.280 ;
        RECT 144.810 156.760 145.455 156.990 ;
        RECT 144.810 155.460 145.010 156.760 ;
        RECT 145.610 155.910 145.810 158.050 ;
        RECT 145.410 155.700 145.810 155.910 ;
        RECT 145.165 155.470 145.810 155.700 ;
        RECT 144.410 155.420 145.010 155.460 ;
        RECT 144.375 154.510 145.010 155.420 ;
        RECT 145.410 155.310 145.810 155.470 ;
        RECT 142.010 153.660 142.410 154.510 ;
        RECT 144.375 154.460 145.310 154.510 ;
        RECT 144.810 154.410 145.310 154.460 ;
        RECT 146.510 154.460 147.210 165.460 ;
        RECT 153.700 162.100 155.400 162.300 ;
        RECT 153.700 160.500 157.100 162.100 ;
        RECT 153.700 160.300 155.400 160.500 ;
        RECT 144.810 154.260 145.455 154.410 ;
        RECT 144.410 154.130 145.810 154.260 ;
        RECT 141.010 153.460 142.410 153.660 ;
        RECT 140.510 153.060 142.410 153.460 ;
        RECT 144.375 153.170 145.810 154.130 ;
        RECT 141.555 152.920 142.365 153.060 ;
        RECT 141.010 152.670 141.410 152.810 ;
        RECT 140.510 152.160 140.810 152.460 ;
        RECT 141.010 152.440 141.845 152.670 ;
        RECT 142.610 152.510 142.910 153.010 ;
        RECT 141.010 152.410 141.410 152.440 ;
        RECT 140.510 151.310 140.710 152.160 ;
        RECT 141.555 152.060 142.365 152.190 ;
        RECT 141.310 151.980 142.710 152.060 ;
        RECT 141.310 151.960 142.840 151.980 ;
        RECT 141.310 151.710 142.910 151.960 ;
        RECT 141.035 151.660 142.910 151.710 ;
        RECT 141.035 151.560 142.710 151.660 ;
        RECT 141.035 151.480 141.845 151.560 ;
        RECT 140.510 150.910 140.810 151.310 ;
        RECT 140.510 150.860 140.710 150.910 ;
        RECT 142.010 150.810 142.410 151.560 ;
        RECT 135.905 150.260 139.010 150.350 ;
        RECT 135.905 150.120 138.465 150.260 ;
        RECT 133.710 149.060 135.010 149.210 ;
        RECT 133.635 148.830 136.195 149.060 ;
        RECT 133.710 148.810 135.010 148.830 ;
        RECT 133.160 147.820 133.390 148.780 ;
        RECT 133.160 146.530 133.390 147.490 ;
        RECT 134.510 146.480 135.010 148.810 ;
        RECT 135.905 147.540 138.465 147.770 ;
        RECT 133.635 146.460 136.195 146.480 ;
        RECT 133.635 146.360 136.210 146.460 ;
        RECT 133.210 146.250 136.210 146.360 ;
        RECT 133.210 146.200 133.910 146.250 ;
        RECT 133.160 145.460 133.910 146.200 ;
        RECT 135.010 145.760 135.310 145.810 ;
        RECT 133.160 145.240 133.390 145.460 ;
        RECT 130.410 142.670 130.710 142.760 ;
        RECT 130.375 141.710 130.710 142.670 ;
        RECT 130.410 141.660 130.710 141.710 ;
        RECT 135.010 141.660 135.410 145.760 ;
        RECT 135.910 145.190 136.210 146.250 ;
        RECT 136.810 145.460 137.310 147.540 ;
        RECT 138.710 146.560 139.010 150.260 ;
        RECT 138.710 146.530 138.940 146.560 ;
        RECT 138.710 146.160 138.940 146.200 ;
        RECT 138.010 145.240 138.940 146.160 ;
        RECT 138.010 145.190 138.910 145.240 ;
        RECT 135.905 145.060 138.910 145.190 ;
        RECT 135.905 144.960 138.465 145.060 ;
        RECT 143.110 143.710 143.510 153.010 ;
        RECT 144.410 152.960 145.810 153.170 ;
        RECT 146.510 153.060 147.110 154.460 ;
        RECT 146.510 153.050 148.110 153.060 ;
        RECT 145.165 152.890 145.725 152.960 ;
        RECT 144.895 152.360 145.455 152.550 ;
        RECT 144.410 152.170 145.610 152.360 ;
        RECT 144.375 151.260 145.610 152.170 ;
        RECT 146.510 151.950 148.900 153.050 ;
        RECT 144.375 151.210 145.725 151.260 ;
        RECT 144.410 151.160 145.725 151.210 ;
        RECT 144.410 151.060 145.810 151.160 ;
        RECT 144.410 150.880 144.910 151.060 ;
        RECT 145.165 151.030 145.810 151.060 ;
        RECT 144.375 150.760 144.910 150.880 ;
        RECT 145.210 150.810 145.810 151.030 ;
        RECT 144.375 149.920 144.610 150.760 ;
        RECT 144.410 149.590 144.610 149.920 ;
        RECT 144.375 148.630 144.610 149.590 ;
        RECT 144.410 148.300 144.610 148.630 ;
        RECT 144.375 147.340 144.610 148.300 ;
        RECT 144.410 147.010 144.610 147.340 ;
        RECT 144.375 146.050 144.610 147.010 ;
        RECT 144.410 145.820 144.610 146.050 ;
        RECT 144.375 144.960 144.610 145.820 ;
        RECT 144.810 149.970 145.410 150.110 ;
        RECT 144.810 149.740 145.455 149.970 ;
        RECT 144.810 149.610 145.410 149.740 ;
        RECT 144.810 147.390 145.010 149.610 ;
        RECT 145.610 148.680 145.810 150.810 ;
        RECT 145.165 148.450 145.810 148.680 ;
        RECT 144.810 147.160 145.455 147.390 ;
        RECT 144.375 144.860 144.605 144.960 ;
        RECT 144.810 144.810 145.010 147.160 ;
        RECT 145.610 146.100 145.810 148.450 ;
        RECT 145.165 145.870 145.810 146.100 ;
        RECT 145.610 145.860 145.810 145.870 ;
        RECT 144.810 144.580 145.455 144.810 ;
        RECT 144.810 144.560 145.410 144.580 ;
        RECT 144.510 144.530 145.410 144.560 ;
        RECT 144.375 144.060 145.410 144.530 ;
        RECT 144.375 143.520 145.710 144.060 ;
        RECT 144.375 143.470 145.725 143.520 ;
        RECT 144.410 143.360 145.725 143.470 ;
        RECT 145.165 143.290 145.725 143.360 ;
        RECT 145.210 143.260 145.710 143.290 ;
        RECT 137.710 142.950 138.610 142.960 ;
        RECT 137.710 142.720 145.725 142.950 ;
        RECT 137.710 141.660 138.610 142.720 ;
        RECT 130.410 141.460 138.610 141.660 ;
        RECT 130.410 141.430 138.455 141.460 ;
        RECT 130.410 141.360 131.710 141.430 ;
        RECT 130.410 139.060 130.710 141.360 ;
        RECT 135.010 139.080 135.410 141.430 ;
        RECT 142.810 140.370 145.610 140.510 ;
        RECT 138.165 140.140 145.725 140.370 ;
        RECT 142.810 140.110 145.610 140.140 ;
        RECT 137.710 139.080 138.610 139.160 ;
        RECT 130.895 139.060 138.610 139.080 ;
        RECT 130.410 138.850 138.610 139.060 ;
        RECT 130.410 138.800 131.710 138.850 ;
        RECT 130.375 138.760 131.710 138.800 ;
        RECT 130.375 137.860 130.710 138.760 ;
        RECT 130.375 137.840 130.605 137.860 ;
        RECT 135.010 136.660 135.410 138.850 ;
        RECT 137.710 137.790 138.610 138.850 ;
        RECT 146.010 137.860 146.310 145.860 ;
        RECT 146.510 139.960 147.110 151.950 ;
        RECT 137.710 137.660 145.725 137.790 ;
        RECT 138.165 137.560 145.725 137.660 ;
        RECT 134.710 135.660 135.710 136.660 ;
        RECT 124.000 131.400 124.900 131.450 ;
        RECT 121.200 124.300 122.200 125.300 ;
        RECT 124.000 124.300 125.000 131.400 ;
        RECT 127.300 125.300 128.300 126.870 ;
        RECT 125.700 124.700 126.700 125.300 ;
        RECT 125.500 124.300 126.700 124.700 ;
        RECT 127.200 124.300 128.300 125.300 ;
        RECT 140.100 124.300 141.100 125.300 ;
        RECT 145.500 124.400 146.500 136.700 ;
        RECT 119.400 118.200 120.200 123.900 ;
        RECT 121.600 119.750 121.900 124.300 ;
        RECT 119.400 117.200 120.400 118.200 ;
        RECT 119.400 116.650 120.200 117.200 ;
        RECT 119.300 115.850 120.200 116.650 ;
        RECT 119.400 109.700 120.200 115.850 ;
        RECT 122.700 111.550 123.000 122.350 ;
        RECT 123.200 113.230 123.680 123.810 ;
        RECT 124.500 123.730 124.800 124.300 ;
        RECT 125.500 124.200 126.400 124.300 ;
        RECT 124.440 123.470 124.860 123.730 ;
        RECT 125.900 123.600 126.400 124.200 ;
        RECT 124.515 122.970 124.745 123.260 ;
        RECT 124.050 121.900 124.400 122.400 ;
        RECT 124.560 121.425 124.700 122.970 ;
        RECT 125.195 122.565 125.425 122.855 ;
        RECT 124.515 121.135 124.745 121.425 ;
        RECT 124.100 120.065 124.400 120.150 ;
        RECT 124.100 119.750 124.405 120.065 ;
        RECT 124.175 119.415 124.405 119.750 ;
        RECT 124.220 116.765 124.360 119.415 ;
        RECT 124.560 117.845 124.700 121.135 ;
        RECT 125.240 120.965 125.380 122.565 ;
        RECT 125.195 120.675 125.425 120.965 ;
        RECT 125.240 117.845 125.380 120.675 ;
        RECT 124.515 117.555 124.745 117.845 ;
        RECT 125.195 117.555 125.425 117.845 ;
        RECT 124.220 116.475 124.720 116.765 ;
        RECT 124.220 116.465 124.405 116.475 ;
        RECT 124.175 116.175 124.405 116.465 ;
        RECT 123.870 114.740 124.230 115.160 ;
        RECT 123.900 112.450 124.200 114.740 ;
        RECT 124.470 113.290 124.730 113.610 ;
        RECT 124.500 112.350 124.700 113.290 ;
        RECT 125.920 113.230 126.400 123.600 ;
        RECT 124.400 111.850 124.800 112.350 ;
        RECT 127.400 111.900 127.950 124.300 ;
        RECT 139.400 124.000 141.500 124.300 ;
        RECT 146.100 124.000 148.100 124.100 ;
        RECT 135.300 123.750 137.300 123.850 ;
        RECT 131.030 123.500 133.135 123.750 ;
        RECT 135.185 123.500 137.300 123.750 ;
        RECT 131.100 122.920 133.000 123.500 ;
        RECT 135.300 123.450 137.300 123.500 ;
        RECT 131.030 122.670 133.135 122.920 ;
        RECT 135.185 122.670 137.290 122.920 ;
        RECT 135.300 122.090 137.200 122.670 ;
        RECT 131.030 121.840 133.135 122.090 ;
        RECT 135.185 121.840 137.290 122.090 ;
        RECT 131.100 121.260 133.000 121.840 ;
        RECT 131.030 121.010 133.135 121.260 ;
        RECT 135.185 121.010 137.290 121.260 ;
        RECT 135.300 120.430 137.200 121.010 ;
        RECT 131.030 120.180 133.135 120.430 ;
        RECT 135.185 120.180 137.290 120.430 ;
        RECT 131.100 119.600 133.000 120.180 ;
        RECT 131.030 119.350 133.135 119.600 ;
        RECT 135.185 119.350 137.290 119.600 ;
        RECT 135.300 118.770 137.200 119.350 ;
        RECT 131.030 118.520 133.135 118.770 ;
        RECT 135.185 118.520 137.290 118.770 ;
        RECT 131.100 117.940 133.000 118.520 ;
        RECT 131.030 117.690 133.135 117.940 ;
        RECT 135.185 117.690 137.290 117.940 ;
        RECT 132.100 114.600 132.600 114.650 ;
        RECT 122.650 111.450 123.000 111.550 ;
        RECT 121.800 111.150 123.000 111.450 ;
        RECT 121.800 111.010 122.700 111.150 ;
        RECT 125.300 111.010 128.200 111.450 ;
        RECT 121.400 110.820 121.600 110.900 ;
        RECT 121.380 110.530 121.610 110.820 ;
        RECT 121.770 110.780 122.770 111.010 ;
        RECT 125.165 110.900 128.200 111.010 ;
        RECT 123.000 110.850 123.200 110.900 ;
        RECT 124.700 110.850 124.900 110.900 ;
        RECT 123.000 110.820 123.300 110.850 ;
        RECT 121.400 110.500 121.600 110.530 ;
        RECT 121.770 110.340 122.770 110.570 ;
        RECT 122.930 110.530 123.300 110.820 ;
        RECT 123.000 110.450 123.300 110.530 ;
        RECT 124.600 110.820 124.900 110.850 ;
        RECT 124.600 110.530 124.960 110.820 ;
        RECT 125.165 110.780 128.165 110.900 ;
        RECT 128.400 110.820 128.700 110.950 ;
        RECT 124.600 110.450 124.900 110.530 ;
        RECT 125.165 110.340 128.165 110.570 ;
        RECT 128.370 110.550 128.700 110.820 ;
        RECT 128.370 110.530 128.600 110.550 ;
        RECT 128.400 110.500 128.600 110.530 ;
        RECT 121.800 110.100 122.700 110.340 ;
        RECT 119.500 109.650 120.100 109.700 ;
        RECT 121.700 109.500 122.700 110.100 ;
        RECT 125.300 110.030 128.100 110.340 ;
        RECT 125.240 109.770 128.160 110.030 ;
        RECT 125.300 109.600 128.100 109.770 ;
        RECT 125.600 109.550 126.000 109.600 ;
        RECT 126.300 109.550 126.700 109.600 ;
        RECT 127.000 109.550 127.400 109.600 ;
        RECT 127.600 109.550 128.000 109.600 ;
        RECT 132.000 78.000 132.600 114.600 ;
        RECT 135.500 114.100 136.700 117.690 ;
        RECT 135.500 114.050 136.600 114.100 ;
        RECT 137.900 110.950 138.400 123.950 ;
        RECT 139.370 123.750 141.500 124.000 ;
        RECT 146.025 123.750 148.130 124.000 ;
        RECT 139.400 123.700 141.500 123.750 ;
        RECT 139.400 123.170 141.400 123.200 ;
        RECT 146.100 123.170 148.100 123.750 ;
        RECT 139.370 122.920 141.475 123.170 ;
        RECT 146.025 122.920 148.130 123.170 ;
        RECT 139.400 122.340 141.400 122.920 ;
        RECT 139.370 122.090 141.475 122.340 ;
        RECT 146.025 122.090 148.130 122.340 ;
        RECT 146.100 121.510 148.100 122.090 ;
        RECT 139.370 121.260 141.475 121.510 ;
        RECT 146.025 121.260 148.130 121.510 ;
        RECT 139.400 120.680 141.400 121.260 ;
        RECT 146.100 121.200 148.100 121.260 ;
        RECT 146.100 120.680 148.100 120.700 ;
        RECT 139.370 120.430 141.475 120.680 ;
        RECT 146.025 120.430 148.130 120.680 ;
        RECT 139.400 120.400 141.400 120.430 ;
        RECT 139.400 119.850 141.400 119.900 ;
        RECT 146.100 119.850 148.100 120.430 ;
        RECT 139.370 119.600 141.475 119.850 ;
        RECT 146.025 119.600 148.130 119.850 ;
        RECT 139.400 119.020 141.400 119.600 ;
        RECT 139.370 118.770 141.475 119.020 ;
        RECT 146.025 118.770 148.130 119.020 ;
        RECT 146.100 118.190 148.100 118.770 ;
        RECT 139.370 117.940 141.475 118.190 ;
        RECT 146.025 117.940 148.130 118.190 ;
        RECT 139.400 116.630 141.400 117.940 ;
        RECT 146.100 117.900 148.100 117.940 ;
        RECT 139.370 116.380 141.475 116.630 ;
        RECT 146.025 116.380 148.130 116.630 ;
        RECT 146.100 115.800 148.100 116.380 ;
        RECT 139.370 115.550 141.475 115.800 ;
        RECT 146.025 115.550 148.130 115.800 ;
        RECT 139.400 114.970 141.400 115.550 ;
        RECT 146.100 115.500 148.100 115.550 ;
        RECT 139.370 114.720 141.475 114.970 ;
        RECT 146.025 114.720 148.130 114.970 ;
        RECT 139.400 114.600 141.400 114.720 ;
        RECT 146.100 114.140 148.100 114.720 ;
        RECT 139.370 113.890 141.475 114.140 ;
        RECT 146.025 113.890 148.130 114.140 ;
        RECT 139.400 113.310 141.400 113.890 ;
        RECT 146.100 113.800 148.100 113.890 ;
        RECT 139.370 113.060 141.475 113.310 ;
        RECT 146.025 113.060 148.130 113.310 ;
        RECT 139.400 113.000 141.400 113.060 ;
        RECT 137.900 110.250 138.500 110.950 ;
        RECT 138.800 110.900 139.200 113.000 ;
        RECT 139.400 112.480 141.400 112.500 ;
        RECT 146.100 112.480 148.100 113.060 ;
        RECT 139.370 112.230 141.475 112.480 ;
        RECT 146.025 112.230 148.130 112.480 ;
        RECT 139.400 111.650 141.400 112.230 ;
        RECT 146.100 112.200 148.100 112.230 ;
        RECT 139.370 111.400 141.475 111.650 ;
        RECT 146.025 111.400 148.130 111.650 ;
        RECT 138.800 110.820 139.600 110.900 ;
        RECT 146.100 110.820 148.100 111.400 ;
        RECT 138.800 110.570 141.475 110.820 ;
        RECT 146.025 110.570 148.130 110.820 ;
        RECT 138.800 110.500 139.600 110.570 ;
        RECT 146.100 110.500 148.100 110.570 ;
        RECT 147.900 110.100 148.800 110.250 ;
        RECT 146.600 109.500 148.800 110.100 ;
        RECT 146.600 109.450 147.000 109.500 ;
        RECT 147.800 109.100 148.800 109.500 ;
        RECT 131.800 76.900 132.900 78.000 ;
        RECT 132.000 74.650 132.600 76.900 ;
      LAYER via ;
        RECT 109.820 194.510 111.320 195.810 ;
        RECT 107.920 174.010 108.420 175.010 ;
        RECT 107.900 171.000 108.600 172.000 ;
        RECT 119.600 194.400 120.200 195.800 ;
        RECT 121.550 193.800 122.450 194.100 ;
        RECT 123.650 193.800 124.550 194.100 ;
        RECT 125.650 193.800 126.650 194.100 ;
        RECT 127.850 193.800 128.750 194.100 ;
        RECT 130.600 193.800 131.000 194.100 ;
        RECT 119.850 192.100 120.350 192.600 ;
        RECT 121.550 192.000 122.450 192.700 ;
        RECT 123.550 192.000 124.550 192.700 ;
        RECT 125.650 192.000 126.650 192.700 ;
        RECT 127.750 192.000 128.750 192.700 ;
        RECT 121.550 190.600 122.450 190.900 ;
        RECT 123.650 190.600 124.550 190.900 ;
        RECT 125.750 190.600 126.650 190.900 ;
        RECT 127.850 190.600 128.750 190.900 ;
        RECT 121.550 190.000 122.350 190.300 ;
        RECT 123.650 190.000 124.450 190.300 ;
        RECT 125.750 190.000 126.550 190.300 ;
        RECT 127.850 190.000 128.650 190.300 ;
        RECT 140.500 194.800 140.900 195.200 ;
        RECT 145.900 194.800 146.400 195.200 ;
        RECT 130.600 192.100 130.900 192.600 ;
        RECT 130.600 190.600 131.000 190.900 ;
        RECT 138.400 192.100 138.700 192.600 ;
        RECT 119.750 188.300 120.450 188.900 ;
        RECT 121.550 188.300 122.250 188.800 ;
        RECT 123.650 188.300 124.350 188.800 ;
        RECT 125.750 188.300 126.450 188.800 ;
        RECT 127.850 188.400 128.550 188.900 ;
        RECT 121.500 186.900 122.400 187.200 ;
        RECT 123.600 186.900 124.500 187.200 ;
        RECT 125.700 186.900 126.600 187.200 ;
        RECT 127.800 186.900 128.700 187.200 ;
        RECT 121.550 186.200 122.450 186.500 ;
        RECT 123.650 186.200 124.550 186.500 ;
        RECT 125.650 186.100 126.650 186.500 ;
        RECT 127.750 186.200 128.750 186.600 ;
        RECT 119.750 184.400 120.450 185.100 ;
        RECT 121.550 184.500 122.350 185.100 ;
        RECT 123.650 184.500 124.450 185.100 ;
        RECT 125.750 184.500 126.550 185.100 ;
        RECT 127.850 184.500 128.650 185.100 ;
        RECT 121.550 183.000 122.450 183.300 ;
        RECT 123.650 183.000 124.550 183.300 ;
        RECT 130.800 190.000 131.200 190.300 ;
        RECT 130.800 186.800 131.200 187.100 ;
        RECT 125.750 183.000 126.650 183.300 ;
        RECT 127.750 183.100 128.650 183.400 ;
        RECT 129.000 183.000 129.300 183.400 ;
        RECT 129.800 183.000 130.200 183.300 ;
        RECT 130.800 183.200 131.200 183.700 ;
        RECT 131.500 186.300 131.800 186.600 ;
        RECT 129.800 181.800 130.200 182.200 ;
        RECT 143.600 188.200 144.200 188.800 ;
        RECT 145.900 188.200 146.400 188.800 ;
        RECT 140.400 184.600 140.900 185.000 ;
        RECT 132.300 183.300 133.300 183.700 ;
        RECT 131.500 181.700 131.800 182.200 ;
        RECT 142.300 184.600 143.400 185.000 ;
        RECT 136.500 183.200 137.100 183.700 ;
        RECT 134.100 179.800 134.600 180.400 ;
        RECT 138.400 183.200 138.700 183.700 ;
        RECT 141.800 183.200 142.100 183.700 ;
        RECT 140.300 181.700 140.800 182.200 ;
        RECT 146.000 176.800 146.800 179.300 ;
        RECT 143.600 176.100 144.200 176.600 ;
        RECT 145.900 176.100 146.400 176.600 ;
        RECT 133.900 174.000 134.900 174.900 ;
        RECT 127.600 171.200 128.400 171.800 ;
        RECT 129.200 169.100 130.000 169.900 ;
        RECT 134.000 169.100 134.800 169.900 ;
        RECT 143.810 164.960 145.010 165.460 ;
        RECT 146.610 165.060 147.210 165.360 ;
        RECT 129.510 161.260 129.910 161.560 ;
        RECT 127.710 156.860 128.310 157.260 ;
        RECT 110.810 155.860 111.110 156.160 ;
        RECT 132.410 155.760 132.810 156.260 ;
        RECT 139.910 161.260 140.210 161.560 ;
        RECT 138.110 156.860 138.510 157.260 ;
        RECT 137.910 155.760 138.410 156.260 ;
        RECT 138.210 154.560 138.710 154.860 ;
        RECT 139.410 154.460 139.710 154.860 ;
        RECT 134.710 152.160 135.010 152.460 ;
        RECT 137.510 152.160 137.810 152.460 ;
        RECT 110.810 148.760 111.110 149.060 ;
        RECT 108.020 130.510 108.520 131.310 ;
        RECT 108.020 127.610 108.420 128.210 ;
        RECT 107.920 125.910 108.520 126.710 ;
        RECT 108.020 124.410 108.520 125.210 ;
        RECT 132.410 148.660 132.810 149.160 ;
        RECT 139.410 152.460 139.710 152.760 ;
        RECT 145.410 155.360 145.810 155.860 ;
        RECT 153.800 160.500 155.200 162.100 ;
        RECT 146.610 155.360 147.110 155.860 ;
        RECT 142.010 154.060 142.410 154.460 ;
        RECT 144.810 154.060 145.310 154.460 ;
        RECT 141.010 152.460 141.410 152.760 ;
        RECT 142.610 152.560 142.910 152.960 ;
        RECT 143.110 152.560 143.510 152.960 ;
        RECT 137.510 150.760 138.410 151.060 ;
        RECT 139.910 150.960 140.210 151.260 ;
        RECT 140.510 150.960 140.810 151.260 ;
        RECT 142.010 150.860 142.410 151.260 ;
        RECT 133.710 148.860 134.910 149.160 ;
        RECT 135.010 145.460 135.310 145.760 ;
        RECT 136.910 145.560 137.210 145.860 ;
        RECT 135.110 143.860 135.410 144.160 ;
        RECT 147.100 152.000 148.900 153.000 ;
        RECT 145.210 150.860 145.610 151.260 ;
        RECT 144.810 149.660 145.410 150.060 ;
        RECT 146.610 149.660 147.110 150.160 ;
        RECT 143.110 143.760 143.510 144.160 ;
        RECT 142.810 140.160 145.610 140.460 ;
        RECT 146.510 140.160 147.010 140.460 ;
        RECT 134.800 135.800 135.600 136.600 ;
        RECT 145.600 135.800 146.400 136.600 ;
        RECT 124.000 130.500 124.900 131.400 ;
        RECT 121.200 124.500 122.100 125.100 ;
        RECT 145.600 127.600 146.400 128.200 ;
        RECT 127.300 126.000 128.300 126.700 ;
        RECT 125.800 124.500 126.500 125.100 ;
        RECT 140.200 124.500 141.000 125.200 ;
        RECT 145.600 124.600 146.400 125.300 ;
        RECT 110.020 117.410 111.220 118.410 ;
        RECT 119.500 123.300 120.200 123.800 ;
        RECT 123.200 123.300 123.600 123.700 ;
        RECT 121.600 119.800 121.900 120.100 ;
        RECT 122.700 122.000 123.000 122.300 ;
        RECT 119.500 117.300 120.100 118.600 ;
        RECT 124.050 121.950 124.400 122.350 ;
        RECT 124.100 119.800 124.400 120.100 ;
        RECT 123.900 112.500 124.200 112.900 ;
        RECT 124.400 111.900 124.800 112.300 ;
        RECT 135.300 123.500 137.300 123.800 ;
        RECT 137.900 123.400 138.400 123.900 ;
        RECT 127.400 111.950 127.950 112.300 ;
        RECT 132.100 114.000 132.600 114.600 ;
        RECT 138.000 117.100 138.400 117.500 ;
        RECT 122.650 111.200 122.950 111.500 ;
        RECT 125.300 111.100 128.200 111.400 ;
        RECT 123.000 110.500 123.300 110.800 ;
        RECT 124.600 110.500 124.900 110.800 ;
        RECT 128.400 110.600 128.700 110.900 ;
        RECT 132.000 110.500 132.600 110.900 ;
        RECT 119.500 109.700 120.100 110.200 ;
        RECT 121.800 109.700 122.500 110.200 ;
        RECT 125.600 109.600 126.000 110.000 ;
        RECT 126.300 109.600 126.700 110.000 ;
        RECT 127.000 109.600 127.400 110.000 ;
        RECT 127.600 109.600 128.000 110.000 ;
        RECT 139.500 117.100 141.300 117.500 ;
        RECT 138.800 112.500 139.100 112.900 ;
        RECT 137.900 110.300 138.500 110.900 ;
        RECT 147.900 109.300 148.800 110.200 ;
        RECT 131.900 77.000 132.800 77.900 ;
      LAYER met2 ;
        RECT 49.100 196.200 50.500 196.250 ;
        RECT 49.100 196.000 112.700 196.200 ;
        RECT 49.100 194.400 120.300 196.000 ;
        RECT 140.450 194.800 146.450 195.200 ;
        RECT 109.620 194.310 120.300 194.400 ;
        RECT 110.730 194.300 120.300 194.310 ;
        RECT 121.450 193.800 131.050 194.100 ;
        RECT 119.750 192.000 128.800 192.700 ;
        RECT 130.550 192.100 138.750 192.600 ;
        RECT 121.450 190.600 131.050 190.900 ;
        RECT 121.450 190.000 131.250 190.300 ;
        RECT 119.700 188.300 128.650 188.900 ;
        RECT 143.550 188.200 146.450 188.800 ;
        RECT 121.450 187.100 122.450 187.200 ;
        RECT 123.550 187.100 124.550 187.200 ;
        RECT 125.650 187.100 126.650 187.200 ;
        RECT 127.750 187.100 128.750 187.200 ;
        RECT 121.450 186.800 131.250 187.100 ;
        RECT 121.150 186.300 131.850 186.600 ;
        RECT 121.500 186.200 122.500 186.300 ;
        RECT 123.600 186.200 124.600 186.300 ;
        RECT 125.600 186.100 126.700 186.300 ;
        RECT 127.700 186.200 128.800 186.300 ;
        RECT 119.700 184.400 128.750 185.100 ;
        RECT 140.350 184.600 143.450 185.000 ;
        RECT 127.700 183.300 128.700 183.400 ;
        RECT 128.950 183.300 129.350 183.400 ;
        RECT 121.250 183.000 130.250 183.300 ;
        RECT 130.750 183.200 142.150 183.700 ;
        RECT 129.750 181.800 140.850 182.200 ;
        RECT 131.350 181.700 140.850 181.800 ;
        RECT 134.050 179.800 143.200 180.400 ;
        RECT 145.950 176.800 146.850 179.300 ;
        RECT 143.550 176.100 146.450 176.600 ;
        RECT 107.870 175.000 112.480 175.010 ;
        RECT 90.250 174.010 135.070 175.000 ;
        RECT 90.250 173.900 108.800 174.010 ;
        RECT 111.230 174.000 135.070 174.010 ;
        RECT 96.400 171.900 108.650 172.000 ;
        RECT 96.400 171.100 128.500 171.900 ;
        RECT 96.400 171.000 108.650 171.100 ;
        RECT 129.100 169.000 134.900 170.000 ;
        RECT 143.760 165.360 147.210 165.460 ;
        RECT 143.760 165.060 147.260 165.360 ;
        RECT 143.760 164.960 147.210 165.060 ;
        RECT 129.460 161.260 140.260 161.560 ;
        RECT 153.750 160.500 155.250 162.100 ;
        RECT 127.660 156.860 138.560 157.260 ;
        RECT 110.710 155.760 138.460 156.260 ;
        RECT 145.360 155.360 147.160 155.860 ;
        RECT 138.160 154.560 139.760 154.860 ;
        RECT 138.210 154.460 139.760 154.560 ;
        RECT 141.960 154.060 145.410 154.460 ;
        RECT 134.610 152.060 137.910 152.560 ;
        RECT 139.360 152.460 141.460 152.760 ;
        RECT 142.560 152.560 143.560 152.960 ;
        RECT 147.050 152.000 148.950 153.000 ;
        RECT 129.260 151.160 130.760 151.760 ;
        RECT 129.260 151.060 138.410 151.160 ;
        RECT 129.260 150.760 138.460 151.060 ;
        RECT 139.810 150.960 140.860 151.260 ;
        RECT 139.810 150.860 140.710 150.960 ;
        RECT 141.960 150.860 145.660 151.260 ;
        RECT 129.260 150.660 138.410 150.760 ;
        RECT 129.260 149.660 130.760 150.660 ;
        RECT 144.810 150.060 147.160 150.160 ;
        RECT 144.760 149.660 147.160 150.060 ;
        RECT 110.710 148.660 135.010 149.160 ;
        RECT 135.010 145.760 137.260 145.860 ;
        RECT 134.960 145.560 137.260 145.760 ;
        RECT 134.960 145.460 137.210 145.560 ;
        RECT 128.310 144.160 129.810 145.160 ;
        RECT 128.310 143.760 143.560 144.160 ;
        RECT 128.310 142.760 129.810 143.760 ;
        RECT 142.610 140.060 147.110 140.560 ;
        RECT 134.700 135.700 146.500 136.700 ;
        RECT 107.920 131.400 112.480 131.410 ;
        RECT 103.200 130.410 125.000 131.400 ;
        RECT 103.200 130.400 108.400 130.410 ;
        RECT 111.300 130.400 125.000 130.410 ;
        RECT 103.200 128.310 108.900 128.400 ;
        RECT 103.200 128.300 112.480 128.310 ;
        RECT 103.200 127.510 146.500 128.300 ;
        RECT 103.200 127.400 108.900 127.510 ;
        RECT 111.300 127.500 146.500 127.510 ;
        RECT 107.870 126.700 112.480 126.710 ;
        RECT 88.000 126.000 128.350 126.700 ;
        RECT 88.000 125.910 128.300 126.000 ;
        RECT 88.000 125.700 108.000 125.910 ;
        RECT 111.300 125.900 128.300 125.910 ;
        RECT 1.000 125.400 2.400 125.450 ;
        RECT 0.950 125.310 108.150 125.400 ;
        RECT 0.950 125.300 112.480 125.310 ;
        RECT 0.950 124.310 126.700 125.300 ;
        RECT 140.100 124.500 146.500 125.400 ;
        RECT 0.950 124.300 108.150 124.310 ;
        RECT 111.300 124.300 126.700 124.310 ;
        RECT 1.000 124.250 2.400 124.300 ;
        RECT 119.450 123.700 123.600 123.800 ;
        RECT 119.450 123.300 123.650 123.700 ;
        RECT 135.200 123.400 138.450 123.900 ;
        RECT 124.000 122.300 124.450 122.350 ;
        RECT 122.650 122.100 124.450 122.300 ;
        RECT 122.650 122.000 123.050 122.100 ;
        RECT 124.000 121.950 124.450 122.100 ;
        RECT 121.550 119.800 124.450 120.100 ;
        RECT 109.620 118.800 112.480 118.810 ;
        RECT 109.620 117.110 120.400 118.800 ;
        RECT 111.250 117.100 120.400 117.110 ;
        RECT 137.800 117.000 141.400 117.500 ;
        RECT 132.000 114.000 136.800 114.600 ;
        RECT 123.850 112.500 139.150 112.900 ;
        RECT 124.350 111.950 128.000 112.300 ;
        RECT 124.350 111.900 124.850 111.950 ;
        RECT 122.600 111.400 123.000 111.500 ;
        RECT 121.800 111.100 128.250 111.400 ;
        RECT 122.950 110.500 124.950 110.800 ;
        RECT 128.350 110.600 132.650 110.900 ;
        RECT 128.400 110.500 132.650 110.600 ;
        RECT 137.850 110.300 138.550 110.900 ;
        RECT 119.450 109.700 123.400 110.200 ;
        RECT 125.300 110.000 147.000 110.100 ;
        RECT 125.300 109.500 147.050 110.000 ;
        RECT 147.850 109.300 148.850 110.200 ;
        RECT 131.800 76.900 132.900 78.000 ;
      LAYER via2 ;
        RECT 49.100 194.500 50.500 196.200 ;
        RECT 146.000 176.800 146.800 179.300 ;
        RECT 90.300 174.000 91.300 174.900 ;
        RECT 96.500 171.100 97.300 171.900 ;
        RECT 153.800 160.500 155.200 162.100 ;
        RECT 147.100 152.000 148.900 153.000 ;
        RECT 129.310 149.660 130.710 151.760 ;
        RECT 128.410 142.860 129.710 145.060 ;
        RECT 103.300 130.500 104.100 131.300 ;
        RECT 103.300 127.500 104.100 128.300 ;
        RECT 88.100 125.800 88.900 126.600 ;
        RECT 1.000 124.300 2.400 125.400 ;
        RECT 137.900 110.300 138.500 110.900 ;
        RECT 119.600 109.700 120.100 110.200 ;
        RECT 147.900 109.300 148.800 110.200 ;
        RECT 131.900 77.000 132.800 77.900 ;
      LAYER met3 ;
        RECT 49.050 194.475 50.550 196.225 ;
        RECT 88.000 125.700 89.000 223.300 ;
        RECT 0.950 124.275 2.450 125.425 ;
        RECT 90.250 4.050 91.350 175.000 ;
        RECT 96.400 4.000 97.400 172.000 ;
        RECT 103.200 130.400 104.200 222.600 ;
        RECT 145.800 179.350 146.800 179.400 ;
        RECT 145.800 176.750 146.825 179.350 ;
        RECT 111.510 151.760 126.910 169.960 ;
        RECT 145.800 160.700 146.800 176.750 ;
        RECT 155.000 162.150 157.200 162.400 ;
        RECT 145.900 160.550 146.800 160.700 ;
        RECT 147.900 153.200 149.100 161.900 ;
        RECT 153.775 160.450 157.200 162.150 ;
        RECT 147.100 153.050 149.100 153.200 ;
        RECT 147.075 151.950 149.100 153.050 ;
        RECT 129.285 151.760 130.735 151.810 ;
        RECT 147.100 151.800 149.100 151.950 ;
        RECT 111.510 149.660 130.810 151.760 ;
        RECT 111.510 138.100 126.910 149.660 ;
        RECT 129.285 149.610 130.735 149.660 ;
        RECT 128.310 142.760 129.810 145.160 ;
        RECT 103.200 16.800 104.200 128.400 ;
        RECT 119.400 108.200 120.200 110.400 ;
        RECT 137.800 110.200 138.600 111.000 ;
        RECT 147.900 110.250 149.100 151.800 ;
        RECT 147.875 109.250 149.100 110.250 ;
        RECT 147.900 109.200 149.100 109.250 ;
        RECT 119.400 80.600 148.660 108.200 ;
        RECT 119.400 76.300 120.200 80.600 ;
        RECT 131.800 76.900 132.900 78.000 ;
        RECT 119.400 73.900 148.660 76.300 ;
        RECT 119.600 48.700 148.660 73.900 ;
        RECT 134.300 4.600 135.300 17.800 ;
        RECT 155.000 7.600 157.200 160.450 ;
      LAYER via3 ;
        RECT 88.100 222.400 88.900 223.100 ;
        RECT 49.100 194.500 50.500 196.200 ;
        RECT 103.300 221.700 104.100 222.500 ;
        RECT 1.000 124.300 2.400 125.400 ;
        RECT 90.300 4.200 91.300 5.100 ;
        RECT 145.900 160.600 146.800 162.200 ;
        RECT 148.000 160.500 149.000 161.800 ;
        RECT 153.800 160.500 155.200 162.100 ;
        RECT 128.410 142.860 129.710 145.060 ;
        RECT 111.650 138.200 126.770 138.520 ;
        RECT 137.900 110.300 138.500 110.900 ;
        RECT 119.700 80.740 120.020 108.060 ;
        RECT 131.900 77.000 132.800 77.900 ;
        RECT 119.700 48.840 120.020 76.160 ;
        RECT 103.300 16.900 104.100 17.700 ;
        RECT 134.400 16.900 135.200 17.700 ;
        RECT 96.500 4.100 97.300 4.900 ;
        RECT 155.200 7.800 157.000 9.600 ;
        RECT 134.400 4.700 135.200 5.500 ;
      LAYER met4 ;
        RECT 88.630 224.100 88.930 224.760 ;
        RECT 88.000 222.300 89.000 224.100 ;
        RECT 154.870 222.600 155.170 224.760 ;
        RECT 103.200 221.600 155.500 222.600 ;
        RECT 50.500 194.495 50.505 196.205 ;
        RECT 111.905 145.060 126.515 169.565 ;
        RECT 150.795 162.300 151.405 162.305 ;
        RECT 145.150 160.400 155.600 162.300 ;
        RECT 128.310 145.060 129.810 145.160 ;
        RECT 111.905 142.860 129.810 145.060 ;
        RECT 111.905 139.955 126.515 142.860 ;
        RECT 128.310 142.760 129.810 142.860 ;
        RECT 111.570 138.120 126.850 138.600 ;
        RECT 0.995 124.295 1.000 125.405 ;
        RECT 119.620 80.660 120.100 108.140 ;
        RECT 136.400 107.805 138.600 112.100 ;
        RECT 121.455 80.995 148.265 107.805 ;
        RECT 131.800 77.200 132.900 78.000 ;
        RECT 119.620 48.760 120.100 76.240 ;
        RECT 131.200 75.905 133.400 77.200 ;
        RECT 121.455 49.095 148.265 75.905 ;
        RECT 103.200 16.800 135.300 17.800 ;
        RECT 90.250 2.650 91.350 5.150 ;
        RECT 96.400 4.000 113.100 5.000 ;
        RECT 90.320 1.000 90.920 2.650 ;
        RECT 112.400 1.000 113.000 4.000 ;
        RECT 134.300 2.500 135.300 5.600 ;
        RECT 155.000 3.600 157.200 9.800 ;
        RECT 134.480 1.000 135.080 2.500 ;
        RECT 156.560 1.000 157.160 3.600 ;
  END
END tt_um_hugodg_temp_sensor
END LIBRARY

